//
// Verilog description for cell conv, 
// Tue Jan 23 11:42:21 2018
//
// Precision RTL Synthesis , 64-bit 2016.1.1.28//


module conv ( clk, rst, image_rsc_addr, image_rsc_re, image_rsc_data_out, 
              image_rsc_triosy_lz, rows_rsc_z, rows_rsc_triosy_lz, cols_rsc_z, 
              cols_rsc_triosy_lz, kernel_rsc_addr, kernel_rsc_re, 
              kernel_rsc_data_out, kernel_rsc_triosy_lz, sortie_rsc_data_in, 
              sortie_rsc_addr, sortie_rsc_re, sortie_rsc_we, sortie_rsc_data_out, 
              sortie_rsc_triosy_lz ) ;

    input clk ;
    input rst ;
    output [15:0]image_rsc_addr ;
    output image_rsc_re ;
    input [31:0]image_rsc_data_out ;
    output image_rsc_triosy_lz ;
    input [31:0]rows_rsc_z ;
    output rows_rsc_triosy_lz ;
    input [31:0]cols_rsc_z ;
    output cols_rsc_triosy_lz ;
    output [8:0]kernel_rsc_addr ;
    output kernel_rsc_re ;
    input [31:0]kernel_rsc_data_out ;
    output kernel_rsc_triosy_lz ;
    output [31:0]sortie_rsc_data_in ;
    output [16:0]sortie_rsc_addr ;
    output sortie_rsc_re ;
    output sortie_rsc_we ;
    input [31:0]sortie_rsc_data_out ;
    output sortie_rsc_triosy_lz ;

    wire [15:0]image_rsc_addr_1_0;
    wire [8:0]kernel_rsc_addr_1_0;
    wire [31:0]sortie_rsc_data_in_1_0;
    wire \sortie_rsc_addr_1_0(2)  , \sortie_rsc_addr_1_0(1)  , 
         \sortie_rsc_addr_1_0(0)  ;
    wire clk_int;
    wire rst_int;
    wire [31:0]rows_rsc_z_int;
    wire [31:0]cols_rsc_z_int;
    wire [31:0]image_rsc_data_out_int;
    wire [31:0]kernel_rsc_data_out_int;
    wire [31:0]sortie_rsc_data_out_int;
    wire \conv_core_inst_fsm_output(10)  , nx14731z1, nx17963z1, nx36106z1, 
         nx37103z1, nx38100z1, nx39097z1, nx40094z1, nx41091z1, nx42088z1, 
         nx46052z1, nx45055z1, nx44058z1, nx43061z1, nx42064z1, nx41067z1, 
         nx40070z1, nx60001z1, nx4461z1, nx14731z2;



    OBUF sortie_rsc_triosy_lz_obuf (.O (sortie_rsc_triosy_lz), .I (
         \conv_core_inst_fsm_output(10)  )) ;
    OBUF sortie_rsc_we_obuf (.O (sortie_rsc_we), .I (nx4461z1)) ;
    OBUF sortie_rsc_re_obuf (.O (sortie_rsc_re), .I (nx60001z1)) ;
    OBUF \sortie_rsc_addr_obuf(0)  (.O (sortie_rsc_addr[0]), .I (
         \sortie_rsc_addr_1_0(0)  )) ;
    OBUF \sortie_rsc_addr_obuf(1)  (.O (sortie_rsc_addr[1]), .I (
         \sortie_rsc_addr_1_0(1)  )) ;
    OBUF \sortie_rsc_addr_obuf(2)  (.O (sortie_rsc_addr[2]), .I (
         \sortie_rsc_addr_1_0(2)  )) ;
    OBUF \sortie_rsc_addr_obuf(3)  (.O (sortie_rsc_addr[3]), .I (nx40070z1)) ;
    OBUF \sortie_rsc_addr_obuf(4)  (.O (sortie_rsc_addr[4]), .I (nx41067z1)) ;
    OBUF \sortie_rsc_addr_obuf(5)  (.O (sortie_rsc_addr[5]), .I (nx42064z1)) ;
    OBUF \sortie_rsc_addr_obuf(6)  (.O (sortie_rsc_addr[6]), .I (nx43061z1)) ;
    OBUF \sortie_rsc_addr_obuf(7)  (.O (sortie_rsc_addr[7]), .I (nx44058z1)) ;
    OBUF \sortie_rsc_addr_obuf(8)  (.O (sortie_rsc_addr[8]), .I (nx45055z1)) ;
    OBUF \sortie_rsc_addr_obuf(9)  (.O (sortie_rsc_addr[9]), .I (nx46052z1)) ;
    OBUF \sortie_rsc_addr_obuf(10)  (.O (sortie_rsc_addr[10]), .I (nx42088z1)) ;
    OBUF \sortie_rsc_addr_obuf(11)  (.O (sortie_rsc_addr[11]), .I (nx41091z1)) ;
    OBUF \sortie_rsc_addr_obuf(12)  (.O (sortie_rsc_addr[12]), .I (nx40094z1)) ;
    OBUF \sortie_rsc_addr_obuf(13)  (.O (sortie_rsc_addr[13]), .I (nx39097z1)) ;
    OBUF \sortie_rsc_addr_obuf(14)  (.O (sortie_rsc_addr[14]), .I (nx38100z1)) ;
    OBUF \sortie_rsc_addr_obuf(15)  (.O (sortie_rsc_addr[15]), .I (nx37103z1)) ;
    OBUF \sortie_rsc_addr_obuf(16)  (.O (sortie_rsc_addr[16]), .I (nx36106z1)) ;
    OBUF \sortie_rsc_data_in_obuf(0)  (.O (sortie_rsc_data_in[0]), .I (
         sortie_rsc_data_in_1_0[0])) ;
    OBUF \sortie_rsc_data_in_obuf(1)  (.O (sortie_rsc_data_in[1]), .I (
         sortie_rsc_data_in_1_0[1])) ;
    OBUF \sortie_rsc_data_in_obuf(2)  (.O (sortie_rsc_data_in[2]), .I (
         sortie_rsc_data_in_1_0[2])) ;
    OBUF \sortie_rsc_data_in_obuf(3)  (.O (sortie_rsc_data_in[3]), .I (
         sortie_rsc_data_in_1_0[3])) ;
    OBUF \sortie_rsc_data_in_obuf(4)  (.O (sortie_rsc_data_in[4]), .I (
         sortie_rsc_data_in_1_0[4])) ;
    OBUF \sortie_rsc_data_in_obuf(5)  (.O (sortie_rsc_data_in[5]), .I (
         sortie_rsc_data_in_1_0[5])) ;
    OBUF \sortie_rsc_data_in_obuf(6)  (.O (sortie_rsc_data_in[6]), .I (
         sortie_rsc_data_in_1_0[6])) ;
    OBUF \sortie_rsc_data_in_obuf(7)  (.O (sortie_rsc_data_in[7]), .I (
         sortie_rsc_data_in_1_0[7])) ;
    OBUF \sortie_rsc_data_in_obuf(8)  (.O (sortie_rsc_data_in[8]), .I (
         sortie_rsc_data_in_1_0[8])) ;
    OBUF \sortie_rsc_data_in_obuf(9)  (.O (sortie_rsc_data_in[9]), .I (
         sortie_rsc_data_in_1_0[9])) ;
    OBUF \sortie_rsc_data_in_obuf(10)  (.O (sortie_rsc_data_in[10]), .I (
         sortie_rsc_data_in_1_0[10])) ;
    OBUF \sortie_rsc_data_in_obuf(11)  (.O (sortie_rsc_data_in[11]), .I (
         sortie_rsc_data_in_1_0[11])) ;
    OBUF \sortie_rsc_data_in_obuf(12)  (.O (sortie_rsc_data_in[12]), .I (
         sortie_rsc_data_in_1_0[12])) ;
    OBUF \sortie_rsc_data_in_obuf(13)  (.O (sortie_rsc_data_in[13]), .I (
         sortie_rsc_data_in_1_0[13])) ;
    OBUF \sortie_rsc_data_in_obuf(14)  (.O (sortie_rsc_data_in[14]), .I (
         sortie_rsc_data_in_1_0[14])) ;
    OBUF \sortie_rsc_data_in_obuf(15)  (.O (sortie_rsc_data_in[15]), .I (
         sortie_rsc_data_in_1_0[15])) ;
    OBUF \sortie_rsc_data_in_obuf(16)  (.O (sortie_rsc_data_in[16]), .I (
         sortie_rsc_data_in_1_0[16])) ;
    OBUF \sortie_rsc_data_in_obuf(17)  (.O (sortie_rsc_data_in[17]), .I (
         sortie_rsc_data_in_1_0[17])) ;
    OBUF \sortie_rsc_data_in_obuf(18)  (.O (sortie_rsc_data_in[18]), .I (
         sortie_rsc_data_in_1_0[18])) ;
    OBUF \sortie_rsc_data_in_obuf(19)  (.O (sortie_rsc_data_in[19]), .I (
         sortie_rsc_data_in_1_0[19])) ;
    OBUF \sortie_rsc_data_in_obuf(20)  (.O (sortie_rsc_data_in[20]), .I (
         sortie_rsc_data_in_1_0[20])) ;
    OBUF \sortie_rsc_data_in_obuf(21)  (.O (sortie_rsc_data_in[21]), .I (
         sortie_rsc_data_in_1_0[21])) ;
    OBUF \sortie_rsc_data_in_obuf(22)  (.O (sortie_rsc_data_in[22]), .I (
         sortie_rsc_data_in_1_0[22])) ;
    OBUF \sortie_rsc_data_in_obuf(23)  (.O (sortie_rsc_data_in[23]), .I (
         sortie_rsc_data_in_1_0[23])) ;
    OBUF \sortie_rsc_data_in_obuf(24)  (.O (sortie_rsc_data_in[24]), .I (
         sortie_rsc_data_in_1_0[24])) ;
    OBUF \sortie_rsc_data_in_obuf(25)  (.O (sortie_rsc_data_in[25]), .I (
         sortie_rsc_data_in_1_0[25])) ;
    OBUF \sortie_rsc_data_in_obuf(26)  (.O (sortie_rsc_data_in[26]), .I (
         sortie_rsc_data_in_1_0[26])) ;
    OBUF \sortie_rsc_data_in_obuf(27)  (.O (sortie_rsc_data_in[27]), .I (
         sortie_rsc_data_in_1_0[27])) ;
    OBUF \sortie_rsc_data_in_obuf(28)  (.O (sortie_rsc_data_in[28]), .I (
         sortie_rsc_data_in_1_0[28])) ;
    OBUF \sortie_rsc_data_in_obuf(29)  (.O (sortie_rsc_data_in[29]), .I (
         sortie_rsc_data_in_1_0[29])) ;
    OBUF \sortie_rsc_data_in_obuf(30)  (.O (sortie_rsc_data_in[30]), .I (
         sortie_rsc_data_in_1_0[30])) ;
    OBUF \sortie_rsc_data_in_obuf(31)  (.O (sortie_rsc_data_in[31]), .I (
         sortie_rsc_data_in_1_0[31])) ;
    OBUF kernel_rsc_triosy_lz_obuf (.O (kernel_rsc_triosy_lz), .I (
         \conv_core_inst_fsm_output(10)  )) ;
    OBUF kernel_rsc_re_obuf (.O (kernel_rsc_re), .I (nx60001z1)) ;
    OBUF \kernel_rsc_addr_obuf(0)  (.O (kernel_rsc_addr[0]), .I (
         kernel_rsc_addr_1_0[0])) ;
    OBUF \kernel_rsc_addr_obuf(1)  (.O (kernel_rsc_addr[1]), .I (
         kernel_rsc_addr_1_0[1])) ;
    OBUF \kernel_rsc_addr_obuf(2)  (.O (kernel_rsc_addr[2]), .I (
         kernel_rsc_addr_1_0[2])) ;
    OBUF \kernel_rsc_addr_obuf(3)  (.O (kernel_rsc_addr[3]), .I (
         kernel_rsc_addr_1_0[3])) ;
    OBUF \kernel_rsc_addr_obuf(4)  (.O (kernel_rsc_addr[4]), .I (
         kernel_rsc_addr_1_0[4])) ;
    OBUF \kernel_rsc_addr_obuf(5)  (.O (kernel_rsc_addr[5]), .I (
         kernel_rsc_addr_1_0[5])) ;
    OBUF \kernel_rsc_addr_obuf(6)  (.O (kernel_rsc_addr[6]), .I (
         kernel_rsc_addr_1_0[6])) ;
    OBUF \kernel_rsc_addr_obuf(7)  (.O (kernel_rsc_addr[7]), .I (
         kernel_rsc_addr_1_0[7])) ;
    OBUF \kernel_rsc_addr_obuf(8)  (.O (kernel_rsc_addr[8]), .I (
         kernel_rsc_addr_1_0[8])) ;
    OBUF cols_rsc_triosy_lz_obuf (.O (cols_rsc_triosy_lz), .I (
         \conv_core_inst_fsm_output(10)  )) ;
    OBUF rows_rsc_triosy_lz_obuf (.O (rows_rsc_triosy_lz), .I (
         \conv_core_inst_fsm_output(10)  )) ;
    OBUF image_rsc_triosy_lz_obuf (.O (image_rsc_triosy_lz), .I (
         \conv_core_inst_fsm_output(10)  )) ;
    OBUF image_rsc_re_obuf (.O (image_rsc_re), .I (nx17963z1)) ;
    OBUF \image_rsc_addr_obuf(0)  (.O (image_rsc_addr[0]), .I (
         image_rsc_addr_1_0[0])) ;
    OBUF \image_rsc_addr_obuf(1)  (.O (image_rsc_addr[1]), .I (
         image_rsc_addr_1_0[1])) ;
    OBUF \image_rsc_addr_obuf(2)  (.O (image_rsc_addr[2]), .I (
         image_rsc_addr_1_0[2])) ;
    OBUF \image_rsc_addr_obuf(3)  (.O (image_rsc_addr[3]), .I (
         image_rsc_addr_1_0[3])) ;
    OBUF \image_rsc_addr_obuf(4)  (.O (image_rsc_addr[4]), .I (
         image_rsc_addr_1_0[4])) ;
    OBUF \image_rsc_addr_obuf(5)  (.O (image_rsc_addr[5]), .I (
         image_rsc_addr_1_0[5])) ;
    OBUF \image_rsc_addr_obuf(6)  (.O (image_rsc_addr[6]), .I (
         image_rsc_addr_1_0[6])) ;
    OBUF \image_rsc_addr_obuf(7)  (.O (image_rsc_addr[7]), .I (
         image_rsc_addr_1_0[7])) ;
    OBUF \image_rsc_addr_obuf(8)  (.O (image_rsc_addr[8]), .I (
         image_rsc_addr_1_0[8])) ;
    OBUF \image_rsc_addr_obuf(9)  (.O (image_rsc_addr[9]), .I (
         image_rsc_addr_1_0[9])) ;
    OBUF \image_rsc_addr_obuf(10)  (.O (image_rsc_addr[10]), .I (
         image_rsc_addr_1_0[10])) ;
    OBUF \image_rsc_addr_obuf(11)  (.O (image_rsc_addr[11]), .I (
         image_rsc_addr_1_0[11])) ;
    OBUF \image_rsc_addr_obuf(12)  (.O (image_rsc_addr[12]), .I (
         image_rsc_addr_1_0[12])) ;
    OBUF \image_rsc_addr_obuf(13)  (.O (image_rsc_addr[13]), .I (
         image_rsc_addr_1_0[13])) ;
    OBUF \image_rsc_addr_obuf(14)  (.O (image_rsc_addr[14]), .I (
         image_rsc_addr_1_0[14])) ;
    OBUF \image_rsc_addr_obuf(15)  (.O (image_rsc_addr[15]), .I (
         image_rsc_addr_1_0[15])) ;
    IBUF \sortie_rsc_data_out_ibuf(0)  (.O (sortie_rsc_data_out_int[0]), .I (
         sortie_rsc_data_out[0])) ;
    IBUF \sortie_rsc_data_out_ibuf(1)  (.O (sortie_rsc_data_out_int[1]), .I (
         sortie_rsc_data_out[1])) ;
    IBUF \sortie_rsc_data_out_ibuf(2)  (.O (sortie_rsc_data_out_int[2]), .I (
         sortie_rsc_data_out[2])) ;
    IBUF \sortie_rsc_data_out_ibuf(3)  (.O (sortie_rsc_data_out_int[3]), .I (
         sortie_rsc_data_out[3])) ;
    IBUF \sortie_rsc_data_out_ibuf(4)  (.O (sortie_rsc_data_out_int[4]), .I (
         sortie_rsc_data_out[4])) ;
    IBUF \sortie_rsc_data_out_ibuf(5)  (.O (sortie_rsc_data_out_int[5]), .I (
         sortie_rsc_data_out[5])) ;
    IBUF \sortie_rsc_data_out_ibuf(6)  (.O (sortie_rsc_data_out_int[6]), .I (
         sortie_rsc_data_out[6])) ;
    IBUF \sortie_rsc_data_out_ibuf(7)  (.O (sortie_rsc_data_out_int[7]), .I (
         sortie_rsc_data_out[7])) ;
    IBUF \sortie_rsc_data_out_ibuf(8)  (.O (sortie_rsc_data_out_int[8]), .I (
         sortie_rsc_data_out[8])) ;
    IBUF \sortie_rsc_data_out_ibuf(9)  (.O (sortie_rsc_data_out_int[9]), .I (
         sortie_rsc_data_out[9])) ;
    IBUF \sortie_rsc_data_out_ibuf(10)  (.O (sortie_rsc_data_out_int[10]), .I (
         sortie_rsc_data_out[10])) ;
    IBUF \sortie_rsc_data_out_ibuf(11)  (.O (sortie_rsc_data_out_int[11]), .I (
         sortie_rsc_data_out[11])) ;
    IBUF \sortie_rsc_data_out_ibuf(12)  (.O (sortie_rsc_data_out_int[12]), .I (
         sortie_rsc_data_out[12])) ;
    IBUF \sortie_rsc_data_out_ibuf(13)  (.O (sortie_rsc_data_out_int[13]), .I (
         sortie_rsc_data_out[13])) ;
    IBUF \sortie_rsc_data_out_ibuf(14)  (.O (sortie_rsc_data_out_int[14]), .I (
         sortie_rsc_data_out[14])) ;
    IBUF \sortie_rsc_data_out_ibuf(15)  (.O (sortie_rsc_data_out_int[15]), .I (
         sortie_rsc_data_out[15])) ;
    IBUF \sortie_rsc_data_out_ibuf(16)  (.O (sortie_rsc_data_out_int[16]), .I (
         sortie_rsc_data_out[16])) ;
    IBUF \sortie_rsc_data_out_ibuf(17)  (.O (sortie_rsc_data_out_int[17]), .I (
         sortie_rsc_data_out[17])) ;
    IBUF \sortie_rsc_data_out_ibuf(18)  (.O (sortie_rsc_data_out_int[18]), .I (
         sortie_rsc_data_out[18])) ;
    IBUF \sortie_rsc_data_out_ibuf(19)  (.O (sortie_rsc_data_out_int[19]), .I (
         sortie_rsc_data_out[19])) ;
    IBUF \sortie_rsc_data_out_ibuf(20)  (.O (sortie_rsc_data_out_int[20]), .I (
         sortie_rsc_data_out[20])) ;
    IBUF \sortie_rsc_data_out_ibuf(21)  (.O (sortie_rsc_data_out_int[21]), .I (
         sortie_rsc_data_out[21])) ;
    IBUF \sortie_rsc_data_out_ibuf(22)  (.O (sortie_rsc_data_out_int[22]), .I (
         sortie_rsc_data_out[22])) ;
    IBUF \sortie_rsc_data_out_ibuf(23)  (.O (sortie_rsc_data_out_int[23]), .I (
         sortie_rsc_data_out[23])) ;
    IBUF \sortie_rsc_data_out_ibuf(24)  (.O (sortie_rsc_data_out_int[24]), .I (
         sortie_rsc_data_out[24])) ;
    IBUF \sortie_rsc_data_out_ibuf(25)  (.O (sortie_rsc_data_out_int[25]), .I (
         sortie_rsc_data_out[25])) ;
    IBUF \sortie_rsc_data_out_ibuf(26)  (.O (sortie_rsc_data_out_int[26]), .I (
         sortie_rsc_data_out[26])) ;
    IBUF \sortie_rsc_data_out_ibuf(27)  (.O (sortie_rsc_data_out_int[27]), .I (
         sortie_rsc_data_out[27])) ;
    IBUF \sortie_rsc_data_out_ibuf(28)  (.O (sortie_rsc_data_out_int[28]), .I (
         sortie_rsc_data_out[28])) ;
    IBUF \sortie_rsc_data_out_ibuf(29)  (.O (sortie_rsc_data_out_int[29]), .I (
         sortie_rsc_data_out[29])) ;
    IBUF \sortie_rsc_data_out_ibuf(30)  (.O (sortie_rsc_data_out_int[30]), .I (
         sortie_rsc_data_out[30])) ;
    IBUF \sortie_rsc_data_out_ibuf(31)  (.O (sortie_rsc_data_out_int[31]), .I (
         sortie_rsc_data_out[31])) ;
    IBUF \kernel_rsc_data_out_ibuf(0)  (.O (kernel_rsc_data_out_int[0]), .I (
         kernel_rsc_data_out[0])) ;
    IBUF \kernel_rsc_data_out_ibuf(1)  (.O (kernel_rsc_data_out_int[1]), .I (
         kernel_rsc_data_out[1])) ;
    IBUF \kernel_rsc_data_out_ibuf(2)  (.O (kernel_rsc_data_out_int[2]), .I (
         kernel_rsc_data_out[2])) ;
    IBUF \kernel_rsc_data_out_ibuf(3)  (.O (kernel_rsc_data_out_int[3]), .I (
         kernel_rsc_data_out[3])) ;
    IBUF \kernel_rsc_data_out_ibuf(4)  (.O (kernel_rsc_data_out_int[4]), .I (
         kernel_rsc_data_out[4])) ;
    IBUF \kernel_rsc_data_out_ibuf(5)  (.O (kernel_rsc_data_out_int[5]), .I (
         kernel_rsc_data_out[5])) ;
    IBUF \kernel_rsc_data_out_ibuf(6)  (.O (kernel_rsc_data_out_int[6]), .I (
         kernel_rsc_data_out[6])) ;
    IBUF \kernel_rsc_data_out_ibuf(7)  (.O (kernel_rsc_data_out_int[7]), .I (
         kernel_rsc_data_out[7])) ;
    IBUF \kernel_rsc_data_out_ibuf(8)  (.O (kernel_rsc_data_out_int[8]), .I (
         kernel_rsc_data_out[8])) ;
    IBUF \kernel_rsc_data_out_ibuf(9)  (.O (kernel_rsc_data_out_int[9]), .I (
         kernel_rsc_data_out[9])) ;
    IBUF \kernel_rsc_data_out_ibuf(10)  (.O (kernel_rsc_data_out_int[10]), .I (
         kernel_rsc_data_out[10])) ;
    IBUF \kernel_rsc_data_out_ibuf(11)  (.O (kernel_rsc_data_out_int[11]), .I (
         kernel_rsc_data_out[11])) ;
    IBUF \kernel_rsc_data_out_ibuf(12)  (.O (kernel_rsc_data_out_int[12]), .I (
         kernel_rsc_data_out[12])) ;
    IBUF \kernel_rsc_data_out_ibuf(13)  (.O (kernel_rsc_data_out_int[13]), .I (
         kernel_rsc_data_out[13])) ;
    IBUF \kernel_rsc_data_out_ibuf(14)  (.O (kernel_rsc_data_out_int[14]), .I (
         kernel_rsc_data_out[14])) ;
    IBUF \kernel_rsc_data_out_ibuf(15)  (.O (kernel_rsc_data_out_int[15]), .I (
         kernel_rsc_data_out[15])) ;
    IBUF \kernel_rsc_data_out_ibuf(16)  (.O (kernel_rsc_data_out_int[16]), .I (
         kernel_rsc_data_out[16])) ;
    IBUF \kernel_rsc_data_out_ibuf(17)  (.O (kernel_rsc_data_out_int[17]), .I (
         kernel_rsc_data_out[17])) ;
    IBUF \kernel_rsc_data_out_ibuf(18)  (.O (kernel_rsc_data_out_int[18]), .I (
         kernel_rsc_data_out[18])) ;
    IBUF \kernel_rsc_data_out_ibuf(19)  (.O (kernel_rsc_data_out_int[19]), .I (
         kernel_rsc_data_out[19])) ;
    IBUF \kernel_rsc_data_out_ibuf(20)  (.O (kernel_rsc_data_out_int[20]), .I (
         kernel_rsc_data_out[20])) ;
    IBUF \kernel_rsc_data_out_ibuf(21)  (.O (kernel_rsc_data_out_int[21]), .I (
         kernel_rsc_data_out[21])) ;
    IBUF \kernel_rsc_data_out_ibuf(22)  (.O (kernel_rsc_data_out_int[22]), .I (
         kernel_rsc_data_out[22])) ;
    IBUF \kernel_rsc_data_out_ibuf(23)  (.O (kernel_rsc_data_out_int[23]), .I (
         kernel_rsc_data_out[23])) ;
    IBUF \kernel_rsc_data_out_ibuf(24)  (.O (kernel_rsc_data_out_int[24]), .I (
         kernel_rsc_data_out[24])) ;
    IBUF \kernel_rsc_data_out_ibuf(25)  (.O (kernel_rsc_data_out_int[25]), .I (
         kernel_rsc_data_out[25])) ;
    IBUF \kernel_rsc_data_out_ibuf(26)  (.O (kernel_rsc_data_out_int[26]), .I (
         kernel_rsc_data_out[26])) ;
    IBUF \kernel_rsc_data_out_ibuf(27)  (.O (kernel_rsc_data_out_int[27]), .I (
         kernel_rsc_data_out[27])) ;
    IBUF \kernel_rsc_data_out_ibuf(28)  (.O (kernel_rsc_data_out_int[28]), .I (
         kernel_rsc_data_out[28])) ;
    IBUF \kernel_rsc_data_out_ibuf(29)  (.O (kernel_rsc_data_out_int[29]), .I (
         kernel_rsc_data_out[29])) ;
    IBUF \kernel_rsc_data_out_ibuf(30)  (.O (kernel_rsc_data_out_int[30]), .I (
         kernel_rsc_data_out[30])) ;
    IBUF \kernel_rsc_data_out_ibuf(31)  (.O (kernel_rsc_data_out_int[31]), .I (
         kernel_rsc_data_out[31])) ;
    IBUF \image_rsc_data_out_ibuf(0)  (.O (image_rsc_data_out_int[0]), .I (
         image_rsc_data_out[0])) ;
    IBUF \image_rsc_data_out_ibuf(1)  (.O (image_rsc_data_out_int[1]), .I (
         image_rsc_data_out[1])) ;
    IBUF \image_rsc_data_out_ibuf(2)  (.O (image_rsc_data_out_int[2]), .I (
         image_rsc_data_out[2])) ;
    IBUF \image_rsc_data_out_ibuf(3)  (.O (image_rsc_data_out_int[3]), .I (
         image_rsc_data_out[3])) ;
    IBUF \image_rsc_data_out_ibuf(4)  (.O (image_rsc_data_out_int[4]), .I (
         image_rsc_data_out[4])) ;
    IBUF \image_rsc_data_out_ibuf(5)  (.O (image_rsc_data_out_int[5]), .I (
         image_rsc_data_out[5])) ;
    IBUF \image_rsc_data_out_ibuf(6)  (.O (image_rsc_data_out_int[6]), .I (
         image_rsc_data_out[6])) ;
    IBUF \image_rsc_data_out_ibuf(7)  (.O (image_rsc_data_out_int[7]), .I (
         image_rsc_data_out[7])) ;
    IBUF \image_rsc_data_out_ibuf(8)  (.O (image_rsc_data_out_int[8]), .I (
         image_rsc_data_out[8])) ;
    IBUF \image_rsc_data_out_ibuf(9)  (.O (image_rsc_data_out_int[9]), .I (
         image_rsc_data_out[9])) ;
    IBUF \image_rsc_data_out_ibuf(10)  (.O (image_rsc_data_out_int[10]), .I (
         image_rsc_data_out[10])) ;
    IBUF \image_rsc_data_out_ibuf(11)  (.O (image_rsc_data_out_int[11]), .I (
         image_rsc_data_out[11])) ;
    IBUF \image_rsc_data_out_ibuf(12)  (.O (image_rsc_data_out_int[12]), .I (
         image_rsc_data_out[12])) ;
    IBUF \image_rsc_data_out_ibuf(13)  (.O (image_rsc_data_out_int[13]), .I (
         image_rsc_data_out[13])) ;
    IBUF \image_rsc_data_out_ibuf(14)  (.O (image_rsc_data_out_int[14]), .I (
         image_rsc_data_out[14])) ;
    IBUF \image_rsc_data_out_ibuf(15)  (.O (image_rsc_data_out_int[15]), .I (
         image_rsc_data_out[15])) ;
    IBUF \image_rsc_data_out_ibuf(16)  (.O (image_rsc_data_out_int[16]), .I (
         image_rsc_data_out[16])) ;
    IBUF \image_rsc_data_out_ibuf(17)  (.O (image_rsc_data_out_int[17]), .I (
         image_rsc_data_out[17])) ;
    IBUF \image_rsc_data_out_ibuf(18)  (.O (image_rsc_data_out_int[18]), .I (
         image_rsc_data_out[18])) ;
    IBUF \image_rsc_data_out_ibuf(19)  (.O (image_rsc_data_out_int[19]), .I (
         image_rsc_data_out[19])) ;
    IBUF \image_rsc_data_out_ibuf(20)  (.O (image_rsc_data_out_int[20]), .I (
         image_rsc_data_out[20])) ;
    IBUF \image_rsc_data_out_ibuf(21)  (.O (image_rsc_data_out_int[21]), .I (
         image_rsc_data_out[21])) ;
    IBUF \image_rsc_data_out_ibuf(22)  (.O (image_rsc_data_out_int[22]), .I (
         image_rsc_data_out[22])) ;
    IBUF \image_rsc_data_out_ibuf(23)  (.O (image_rsc_data_out_int[23]), .I (
         image_rsc_data_out[23])) ;
    IBUF \image_rsc_data_out_ibuf(24)  (.O (image_rsc_data_out_int[24]), .I (
         image_rsc_data_out[24])) ;
    IBUF \image_rsc_data_out_ibuf(25)  (.O (image_rsc_data_out_int[25]), .I (
         image_rsc_data_out[25])) ;
    IBUF \image_rsc_data_out_ibuf(26)  (.O (image_rsc_data_out_int[26]), .I (
         image_rsc_data_out[26])) ;
    IBUF \image_rsc_data_out_ibuf(27)  (.O (image_rsc_data_out_int[27]), .I (
         image_rsc_data_out[27])) ;
    IBUF \image_rsc_data_out_ibuf(28)  (.O (image_rsc_data_out_int[28]), .I (
         image_rsc_data_out[28])) ;
    IBUF \image_rsc_data_out_ibuf(29)  (.O (image_rsc_data_out_int[29]), .I (
         image_rsc_data_out[29])) ;
    IBUF \image_rsc_data_out_ibuf(30)  (.O (image_rsc_data_out_int[30]), .I (
         image_rsc_data_out[30])) ;
    IBUF \image_rsc_data_out_ibuf(31)  (.O (image_rsc_data_out_int[31]), .I (
         image_rsc_data_out[31])) ;
    IBUF \cols_rsc_z_ibuf(0)  (.O (cols_rsc_z_int[0]), .I (cols_rsc_z[0])) ;
    IBUF \cols_rsc_z_ibuf(1)  (.O (cols_rsc_z_int[1]), .I (cols_rsc_z[1])) ;
    IBUF \cols_rsc_z_ibuf(2)  (.O (cols_rsc_z_int[2]), .I (cols_rsc_z[2])) ;
    IBUF \cols_rsc_z_ibuf(3)  (.O (cols_rsc_z_int[3]), .I (cols_rsc_z[3])) ;
    IBUF \cols_rsc_z_ibuf(4)  (.O (cols_rsc_z_int[4]), .I (cols_rsc_z[4])) ;
    IBUF \cols_rsc_z_ibuf(5)  (.O (cols_rsc_z_int[5]), .I (cols_rsc_z[5])) ;
    IBUF \cols_rsc_z_ibuf(6)  (.O (cols_rsc_z_int[6]), .I (cols_rsc_z[6])) ;
    IBUF \cols_rsc_z_ibuf(7)  (.O (cols_rsc_z_int[7]), .I (cols_rsc_z[7])) ;
    IBUF \cols_rsc_z_ibuf(8)  (.O (cols_rsc_z_int[8]), .I (cols_rsc_z[8])) ;
    IBUF \cols_rsc_z_ibuf(9)  (.O (cols_rsc_z_int[9]), .I (cols_rsc_z[9])) ;
    IBUF \cols_rsc_z_ibuf(10)  (.O (cols_rsc_z_int[10]), .I (cols_rsc_z[10])) ;
    IBUF \cols_rsc_z_ibuf(11)  (.O (cols_rsc_z_int[11]), .I (cols_rsc_z[11])) ;
    IBUF \cols_rsc_z_ibuf(12)  (.O (cols_rsc_z_int[12]), .I (cols_rsc_z[12])) ;
    IBUF \cols_rsc_z_ibuf(13)  (.O (cols_rsc_z_int[13]), .I (cols_rsc_z[13])) ;
    IBUF \cols_rsc_z_ibuf(14)  (.O (cols_rsc_z_int[14]), .I (cols_rsc_z[14])) ;
    IBUF \cols_rsc_z_ibuf(15)  (.O (cols_rsc_z_int[15]), .I (cols_rsc_z[15])) ;
    IBUF \cols_rsc_z_ibuf(16)  (.O (cols_rsc_z_int[16]), .I (cols_rsc_z[16])) ;
    IBUF \cols_rsc_z_ibuf(17)  (.O (cols_rsc_z_int[17]), .I (cols_rsc_z[17])) ;
    IBUF \cols_rsc_z_ibuf(18)  (.O (cols_rsc_z_int[18]), .I (cols_rsc_z[18])) ;
    IBUF \cols_rsc_z_ibuf(19)  (.O (cols_rsc_z_int[19]), .I (cols_rsc_z[19])) ;
    IBUF \cols_rsc_z_ibuf(20)  (.O (cols_rsc_z_int[20]), .I (cols_rsc_z[20])) ;
    IBUF \cols_rsc_z_ibuf(21)  (.O (cols_rsc_z_int[21]), .I (cols_rsc_z[21])) ;
    IBUF \cols_rsc_z_ibuf(22)  (.O (cols_rsc_z_int[22]), .I (cols_rsc_z[22])) ;
    IBUF \cols_rsc_z_ibuf(23)  (.O (cols_rsc_z_int[23]), .I (cols_rsc_z[23])) ;
    IBUF \cols_rsc_z_ibuf(24)  (.O (cols_rsc_z_int[24]), .I (cols_rsc_z[24])) ;
    IBUF \cols_rsc_z_ibuf(25)  (.O (cols_rsc_z_int[25]), .I (cols_rsc_z[25])) ;
    IBUF \cols_rsc_z_ibuf(26)  (.O (cols_rsc_z_int[26]), .I (cols_rsc_z[26])) ;
    IBUF \cols_rsc_z_ibuf(27)  (.O (cols_rsc_z_int[27]), .I (cols_rsc_z[27])) ;
    IBUF \cols_rsc_z_ibuf(28)  (.O (cols_rsc_z_int[28]), .I (cols_rsc_z[28])) ;
    IBUF \cols_rsc_z_ibuf(29)  (.O (cols_rsc_z_int[29]), .I (cols_rsc_z[29])) ;
    IBUF \cols_rsc_z_ibuf(30)  (.O (cols_rsc_z_int[30]), .I (cols_rsc_z[30])) ;
    IBUF \cols_rsc_z_ibuf(31)  (.O (cols_rsc_z_int[31]), .I (cols_rsc_z[31])) ;
    IBUF \rows_rsc_z_ibuf(0)  (.O (rows_rsc_z_int[0]), .I (rows_rsc_z[0])) ;
    IBUF \rows_rsc_z_ibuf(1)  (.O (rows_rsc_z_int[1]), .I (rows_rsc_z[1])) ;
    IBUF \rows_rsc_z_ibuf(2)  (.O (rows_rsc_z_int[2]), .I (rows_rsc_z[2])) ;
    IBUF \rows_rsc_z_ibuf(3)  (.O (rows_rsc_z_int[3]), .I (rows_rsc_z[3])) ;
    IBUF \rows_rsc_z_ibuf(4)  (.O (rows_rsc_z_int[4]), .I (rows_rsc_z[4])) ;
    IBUF \rows_rsc_z_ibuf(5)  (.O (rows_rsc_z_int[5]), .I (rows_rsc_z[5])) ;
    IBUF \rows_rsc_z_ibuf(6)  (.O (rows_rsc_z_int[6]), .I (rows_rsc_z[6])) ;
    IBUF \rows_rsc_z_ibuf(7)  (.O (rows_rsc_z_int[7]), .I (rows_rsc_z[7])) ;
    IBUF \rows_rsc_z_ibuf(8)  (.O (rows_rsc_z_int[8]), .I (rows_rsc_z[8])) ;
    IBUF \rows_rsc_z_ibuf(9)  (.O (rows_rsc_z_int[9]), .I (rows_rsc_z[9])) ;
    IBUF \rows_rsc_z_ibuf(10)  (.O (rows_rsc_z_int[10]), .I (rows_rsc_z[10])) ;
    IBUF \rows_rsc_z_ibuf(11)  (.O (rows_rsc_z_int[11]), .I (rows_rsc_z[11])) ;
    IBUF \rows_rsc_z_ibuf(12)  (.O (rows_rsc_z_int[12]), .I (rows_rsc_z[12])) ;
    IBUF \rows_rsc_z_ibuf(13)  (.O (rows_rsc_z_int[13]), .I (rows_rsc_z[13])) ;
    IBUF \rows_rsc_z_ibuf(14)  (.O (rows_rsc_z_int[14]), .I (rows_rsc_z[14])) ;
    IBUF \rows_rsc_z_ibuf(15)  (.O (rows_rsc_z_int[15]), .I (rows_rsc_z[15])) ;
    IBUF \rows_rsc_z_ibuf(16)  (.O (rows_rsc_z_int[16]), .I (rows_rsc_z[16])) ;
    IBUF \rows_rsc_z_ibuf(17)  (.O (rows_rsc_z_int[17]), .I (rows_rsc_z[17])) ;
    IBUF \rows_rsc_z_ibuf(18)  (.O (rows_rsc_z_int[18]), .I (rows_rsc_z[18])) ;
    IBUF \rows_rsc_z_ibuf(19)  (.O (rows_rsc_z_int[19]), .I (rows_rsc_z[19])) ;
    IBUF \rows_rsc_z_ibuf(20)  (.O (rows_rsc_z_int[20]), .I (rows_rsc_z[20])) ;
    IBUF \rows_rsc_z_ibuf(21)  (.O (rows_rsc_z_int[21]), .I (rows_rsc_z[21])) ;
    IBUF \rows_rsc_z_ibuf(22)  (.O (rows_rsc_z_int[22]), .I (rows_rsc_z[22])) ;
    IBUF \rows_rsc_z_ibuf(23)  (.O (rows_rsc_z_int[23]), .I (rows_rsc_z[23])) ;
    IBUF \rows_rsc_z_ibuf(24)  (.O (rows_rsc_z_int[24]), .I (rows_rsc_z[24])) ;
    IBUF \rows_rsc_z_ibuf(25)  (.O (rows_rsc_z_int[25]), .I (rows_rsc_z[25])) ;
    IBUF \rows_rsc_z_ibuf(26)  (.O (rows_rsc_z_int[26]), .I (rows_rsc_z[26])) ;
    IBUF \rows_rsc_z_ibuf(27)  (.O (rows_rsc_z_int[27]), .I (rows_rsc_z[27])) ;
    IBUF \rows_rsc_z_ibuf(28)  (.O (rows_rsc_z_int[28]), .I (rows_rsc_z[28])) ;
    IBUF \rows_rsc_z_ibuf(29)  (.O (rows_rsc_z_int[29]), .I (rows_rsc_z[29])) ;
    IBUF \rows_rsc_z_ibuf(30)  (.O (rows_rsc_z_int[30]), .I (rows_rsc_z[30])) ;
    IBUF \rows_rsc_z_ibuf(31)  (.O (rows_rsc_z_int[31]), .I (rows_rsc_z[31])) ;
    IBUF rst_ibuf (.O (rst_int), .I (rst)) ;
    GND ps_gnd (.G (nx14731z1)) ;
    VCC ps_vcc (.P (nx14731z2)) ;
    conv_core_0 conv_core_inst (.px1550 (nx4461z1), .px1549 (nx60001z1), .px1548 (
                nx40070z1), .px1547 (nx41067z1), .px1546 (nx42064z1), .px1545 (
                nx43061z1), .px1544 (nx44058z1), .px1543 (nx45055z1), .px1542 (
                nx46052z1), .px1541 (nx42088z1), .px1540 (nx41091z1), .px1539 (
                nx40094z1), .px1538 (nx39097z1), .px1537 (nx38100z1), .px1536 (
                nx37103z1), .px1535 (nx36106z1), .px1534 (nx17963z1), .p_nbus_image_rsc_data_out_int (
                {image_rsc_data_out_int[16],image_rsc_data_out_int[15],
                image_rsc_data_out_int[14],image_rsc_data_out_int[13],
                image_rsc_data_out_int[12],image_rsc_data_out_int[11],
                image_rsc_data_out_int[10],image_rsc_data_out_int[9],
                image_rsc_data_out_int[8],image_rsc_data_out_int[7],
                image_rsc_data_out_int[6],image_rsc_data_out_int[5],
                image_rsc_data_out_int[4],image_rsc_data_out_int[3],
                image_rsc_data_out_int[2],image_rsc_data_out_int[1],
                image_rsc_data_out_int[0],image_rsc_data_out_int[31],
                image_rsc_data_out_int[30],image_rsc_data_out_int[29],
                image_rsc_data_out_int[28],image_rsc_data_out_int[27],
                image_rsc_data_out_int[26],image_rsc_data_out_int[25],
                image_rsc_data_out_int[24],image_rsc_data_out_int[23],
                image_rsc_data_out_int[22],image_rsc_data_out_int[21],
                image_rsc_data_out_int[20],image_rsc_data_out_int[19],
                image_rsc_data_out_int[18],image_rsc_data_out_int[17]}), .\p_fsm_output(10)   (
                \conv_core_inst_fsm_output(10)  ), .\p_sortie_rsc_addr_1_0(0)   (
                \sortie_rsc_addr_1_0(0)  ), .\p_sortie_rsc_addr_1_0(1)   (
                \sortie_rsc_addr_1_0(1)  ), .\p_sortie_rsc_addr_1_0(2)   (
                \sortie_rsc_addr_1_0(2)  ), .p_nbus_cols_rsc_z_int ({
                cols_rsc_z_int[0],cols_rsc_z_int[1],cols_rsc_z_int[2],
                cols_rsc_z_int[3],cols_rsc_z_int[4],cols_rsc_z_int[5],
                cols_rsc_z_int[6],cols_rsc_z_int[7],cols_rsc_z_int[8],
                cols_rsc_z_int[9],cols_rsc_z_int[10],cols_rsc_z_int[11],
                cols_rsc_z_int[12],cols_rsc_z_int[13],cols_rsc_z_int[14],
                cols_rsc_z_int[15],cols_rsc_z_int[16],cols_rsc_z_int[17],
                cols_rsc_z_int[18],cols_rsc_z_int[19],cols_rsc_z_int[20],
                cols_rsc_z_int[21],cols_rsc_z_int[22],cols_rsc_z_int[23],
                cols_rsc_z_int[24],cols_rsc_z_int[25],cols_rsc_z_int[26],
                cols_rsc_z_int[27],cols_rsc_z_int[28],cols_rsc_z_int[29],
                cols_rsc_z_int[30],cols_rsc_z_int[31]}), .p_nbus_rows_rsc_z_int (
                {rows_rsc_z_int[0],rows_rsc_z_int[1],rows_rsc_z_int[2],
                rows_rsc_z_int[3],rows_rsc_z_int[4],rows_rsc_z_int[5],
                rows_rsc_z_int[6],rows_rsc_z_int[7],rows_rsc_z_int[8],
                rows_rsc_z_int[9],rows_rsc_z_int[10],rows_rsc_z_int[11],
                rows_rsc_z_int[12],rows_rsc_z_int[13],rows_rsc_z_int[14],
                rows_rsc_z_int[15],rows_rsc_z_int[16],rows_rsc_z_int[17],
                rows_rsc_z_int[18],rows_rsc_z_int[19],rows_rsc_z_int[20],
                rows_rsc_z_int[21],rows_rsc_z_int[22],rows_rsc_z_int[23],
                rows_rsc_z_int[24],rows_rsc_z_int[25],rows_rsc_z_int[26],
                rows_rsc_z_int[27],rows_rsc_z_int[28],rows_rsc_z_int[29],
                rows_rsc_z_int[30],rows_rsc_z_int[31]}), .p_nbus_image_rsc_addr_1_0 (
                {image_rsc_addr_1_0[0],image_rsc_addr_1_0[1],
                image_rsc_addr_1_0[2],image_rsc_addr_1_0[15],
                image_rsc_addr_1_0[14],image_rsc_addr_1_0[13],
                image_rsc_addr_1_0[12],image_rsc_addr_1_0[11],
                image_rsc_addr_1_0[10],image_rsc_addr_1_0[9],
                image_rsc_addr_1_0[8],image_rsc_addr_1_0[7],
                image_rsc_addr_1_0[6],image_rsc_addr_1_0[5],
                image_rsc_addr_1_0[4],image_rsc_addr_1_0[3]}), .p_nbus_kernel_rsc_data_out_int (
                {kernel_rsc_data_out_int[0],kernel_rsc_data_out_int[1],
                kernel_rsc_data_out_int[2],kernel_rsc_data_out_int[3],
                kernel_rsc_data_out_int[4],kernel_rsc_data_out_int[5],
                kernel_rsc_data_out_int[6],kernel_rsc_data_out_int[7],
                kernel_rsc_data_out_int[8],kernel_rsc_data_out_int[9],
                kernel_rsc_data_out_int[10],kernel_rsc_data_out_int[11],
                kernel_rsc_data_out_int[12],kernel_rsc_data_out_int[13],
                kernel_rsc_data_out_int[14],kernel_rsc_data_out_int[15],
                kernel_rsc_data_out_int[16],kernel_rsc_data_out_int[17],
                kernel_rsc_data_out_int[18],kernel_rsc_data_out_int[19],
                kernel_rsc_data_out_int[20],kernel_rsc_data_out_int[21],
                kernel_rsc_data_out_int[22],kernel_rsc_data_out_int[23],
                kernel_rsc_data_out_int[24],kernel_rsc_data_out_int[25],
                kernel_rsc_data_out_int[26],kernel_rsc_data_out_int[27],
                kernel_rsc_data_out_int[28],kernel_rsc_data_out_int[29],
                kernel_rsc_data_out_int[30],kernel_rsc_data_out_int[31]}), .p_nbus_sortie_rsc_data_out_int (
                {sortie_rsc_data_out_int[0],sortie_rsc_data_out_int[1],
                sortie_rsc_data_out_int[2],sortie_rsc_data_out_int[3],
                sortie_rsc_data_out_int[4],sortie_rsc_data_out_int[5],
                sortie_rsc_data_out_int[6],sortie_rsc_data_out_int[7],
                sortie_rsc_data_out_int[8],sortie_rsc_data_out_int[9],
                sortie_rsc_data_out_int[10],sortie_rsc_data_out_int[11],
                sortie_rsc_data_out_int[12],sortie_rsc_data_out_int[13],
                sortie_rsc_data_out_int[14],sortie_rsc_data_out_int[15],
                sortie_rsc_data_out_int[16],sortie_rsc_data_out_int[17],
                sortie_rsc_data_out_int[18],sortie_rsc_data_out_int[19],
                sortie_rsc_data_out_int[20],sortie_rsc_data_out_int[21],
                sortie_rsc_data_out_int[22],sortie_rsc_data_out_int[23],
                sortie_rsc_data_out_int[24],sortie_rsc_data_out_int[25],
                sortie_rsc_data_out_int[26],sortie_rsc_data_out_int[27],
                sortie_rsc_data_out_int[28],sortie_rsc_data_out_int[29],
                sortie_rsc_data_out_int[30],sortie_rsc_data_out_int[31]}), .p_rst_int (
                rst_int), .p_clk_int (clk_int), .p_nbus_sortie_rsc_data_in_1_0 (
                {sortie_rsc_data_in_1_0[31],sortie_rsc_data_in_1_0[30],
                sortie_rsc_data_in_1_0[29],sortie_rsc_data_in_1_0[28],
                sortie_rsc_data_in_1_0[27],sortie_rsc_data_in_1_0[26],
                sortie_rsc_data_in_1_0[25],sortie_rsc_data_in_1_0[24],
                sortie_rsc_data_in_1_0[23],sortie_rsc_data_in_1_0[22],
                sortie_rsc_data_in_1_0[21],sortie_rsc_data_in_1_0[20],
                sortie_rsc_data_in_1_0[19],sortie_rsc_data_in_1_0[18],
                sortie_rsc_data_in_1_0[17],sortie_rsc_data_in_1_0[16],
                sortie_rsc_data_in_1_0[15],sortie_rsc_data_in_1_0[14],
                sortie_rsc_data_in_1_0[13],sortie_rsc_data_in_1_0[12],
                sortie_rsc_data_in_1_0[11],sortie_rsc_data_in_1_0[10],
                sortie_rsc_data_in_1_0[9],sortie_rsc_data_in_1_0[8],
                sortie_rsc_data_in_1_0[7],sortie_rsc_data_in_1_0[6],
                sortie_rsc_data_in_1_0[5],sortie_rsc_data_in_1_0[4],
                sortie_rsc_data_in_1_0[3],sortie_rsc_data_in_1_0[2],
                sortie_rsc_data_in_1_0[1],sortie_rsc_data_in_1_0[0]}), .p_nbus_kernel_rsc_addr_1_0 (
                {kernel_rsc_addr_1_0[8],kernel_rsc_addr_1_0[7],
                kernel_rsc_addr_1_0[6],kernel_rsc_addr_1_0[5],
                kernel_rsc_addr_1_0[4],kernel_rsc_addr_1_0[3],
                kernel_rsc_addr_1_0[2],kernel_rsc_addr_1_0[1],
                kernel_rsc_addr_1_0[0]}), .px1140 (nx14731z1), .px1551 (
                nx14731z2)) ;
    BUFGP clk_ibuf (.O (clk_int), .I (clk)) ;
endmodule


module conv_core_0 ( px1550, px1549, px1548, px1547, px1546, px1545, px1544, 
                     px1543, px1542, px1541, px1540, px1539, px1538, px1537, 
                     px1536, px1535, px1534, p_nbus_image_rsc_data_out_int, 
                     \p_fsm_output(10)  , \p_sortie_rsc_addr_1_0(0)  , 
                     \p_sortie_rsc_addr_1_0(1)  , \p_sortie_rsc_addr_1_0(2)  , 
                     p_nbus_cols_rsc_z_int, p_nbus_rows_rsc_z_int, 
                     p_nbus_image_rsc_addr_1_0, p_nbus_kernel_rsc_data_out_int, 
                     p_nbus_sortie_rsc_data_out_int, p_rst_int, p_clk_int, 
                     p_nbus_sortie_rsc_data_in_1_0, p_nbus_kernel_rsc_addr_1_0, 
                     px1140, px1551 ) ;

    output px1550 ;
    output px1549 ;
    output px1548 ;
    output px1547 ;
    output px1546 ;
    output px1545 ;
    output px1544 ;
    output px1543 ;
    output px1542 ;
    output px1541 ;
    output px1540 ;
    output px1539 ;
    output px1538 ;
    output px1537 ;
    output px1536 ;
    output px1535 ;
    output px1534 ;
    input [31:0]p_nbus_image_rsc_data_out_int ;
    output \p_fsm_output(10)   ;
    output \p_sortie_rsc_addr_1_0(0)   ;
    output \p_sortie_rsc_addr_1_0(1)   ;
    output \p_sortie_rsc_addr_1_0(2)   ;
    input [31:0]p_nbus_cols_rsc_z_int ;
    input [31:0]p_nbus_rows_rsc_z_int ;
    output [15:0]p_nbus_image_rsc_addr_1_0 ;
    input [31:0]p_nbus_kernel_rsc_data_out_int ;
    input [31:0]p_nbus_sortie_rsc_data_out_int ;
    input p_rst_int ;
    input p_clk_int ;
    output [31:0]p_nbus_sortie_rsc_data_in_1_0 ;
    output [8:0]p_nbus_kernel_rsc_addr_1_0 ;
    input px1140 ;
    input px1551 ;

    wire nx6185z1, nx6185z2, nx6185z3, nx6185z4, nx6185z5, nx6185z6, nx6185z7, 
         nx6185z8, nx6185z9, nx6185z10, nx6185z11, nx6185z12, nx6185z13, 
         nx6185z14, nx6185z15, nx6185z16, nx6185z17, nx6185z18, nx6185z19, 
         nx6185z20, nx6185z21, nx6185z22, nx6185z23, nx6185z24, nx6185z25, 
         nx6185z26, nx6185z27, nx6185z28, nx6185z29, nx6185z30, nx6185z31, 
         nx28350z2, nx14411z2, nx13414z2, nx22387z2, nx20393z5, nx18544z3, 
         nx20393z4, nx49642z6, nx49642z3, nx49642z5, nx49641z5, nx49641z4, 
         nx48653z5, nx48653z4, nx48652z5, nx48652z4, nx48651z6, nx48651z5, 
         nx48650z5, nx48650z4, nx48649z5, nx48649z4, nx48648z5, nx48648z4, 
         nx48647z5, nx48647z4, nx48646z5, nx48646z4, nx48645z5, nx48645z4, 
         nx48644z5, nx48644z4, nx47656z5, nx47656z4, nx47655z5, nx47655z4, 
         nx47654z6, nx47654z5, nx47653z5, nx47653z4, nx47652z5, nx47652z4, 
         nx47651z5, nx47651z4, nx47650z5, nx47650z4, nx47649z5, nx47649z4, 
         nx47648z5, nx47648z4, nx47647z5, nx47647z4, nx28341z5, nx28341z4, 
         nx28342z5, nx28342z4, nx28343z5, nx28343z4, nx28344z5, nx28344z4, 
         nx28345z5, nx28345z4, nx28346z5, nx28346z4, nx28347z5, nx28347z4, 
         nx28348z5, nx28348z4, nx28349z5, nx28349z4, nx28350z5, nx28350z4, 
         nx39517z4, nx58321z1, nx39517z6, nx57324z1, nx56327z1, nx55330z1, 
         nx59318z1, nx39520z4, nx21003z2, nx22000z1, nx22997z1, nx23994z1, 
         nx18544z2, nx24991z1, nx21003z1, nx20393z3, nx13414z1, \fsm_output(1)  , 
         nx14411z1, \conv_core_core_fsm_inst_fsm_output(2)  , nx15408z1, 
         \fsm_output(4)  , \fsm_output(5)  , \fsm_output(6)  , nx19396z1, 
         \fsm_output(7)  , nx20393z1, \fsm_output(8)  , nx21390z1, 
         \fsm_output(9)  , nx22387z1, nx43133z1, \fsm_output(0)  , nx12614z2;
    wire [4:0]conv_core_inst_for_for_for_for_n_4_0_sva_3;
    wire nx20538z1, nx19541z1, nx18544z1, nx20393z2, nx60570z1, 
         for_for_for_for_if_for_for_for_for_if_and_2_itm, nx12614z1;
    wire \fsm_output(3)  ;
    wire for_for_for_for_slc_for_for_for_for_acc_5_itm;
    wire [13:0]conv_core_inst_for_for_for_for_if_acc_psp_sva_1;
    wire not_fsm_output_4, nx33183z1, nx32186z1, nx31189z1, nx30192z1, 
         \for_for_j_sva(3)  , nx29195z1, nx28198z1, nx27201z1, nx26204z1, 
         nx25207z1, nx24210z1, nx30218z1, nx31215z1, nx32212z1, nx33209z1, 
         nx34206z1, nx35203z1, nx36200z1, nx37197z1, nx38194z1, nx39191z1, 
         nx41187z1, nx42184z1, nx43181z1, nx44178z1, nx45175z1, nx46172z1, 
         nx47169z1, nx48166z1, nx49163z1, nx50160z1, nx52156z2, nx53153z1, 
         nx52156z1, \for_for_j_sva(31)  ;
    wire [31:0]conv_core_inst_cols_1_sva_1;
    wire nx51642z1;
    wire [31:0]conv_core_inst_for_i_sva;
    wire nx50645z1, nx49648z1, nx48651z1, nx47654z1, nx46657z1, nx45660z1, 
         nx44663z1, nx43666z1, nx42669z1, nx42211z1, nx43208z1, nx44205z1, 
         nx45202z1, nx46199z1, nx47196z1, nx48193z1, nx49190z1, nx50187z1, 
         nx51184z1, nx53180z1, nx54177z1, nx55174z1, nx56171z1, nx57168z1, 
         nx58165z1, nx59162z1, nx60159z1, nx61156z1, nx62153z1, nx64149z2, 
         nx65146z1, nx64149z1;
    wire [31:0]conv_core_inst_rows_1_sva_2;
    wire nx9631z1, nx5701z1, nx4704z1, nx3707z1, nx2710z1;
    wire [4:4]conv_core_inst_for_for_for_for_n_4_0_sva;
    wire nx1713z1, \for_for_for_for_n_4_0_sva(4)  ;
    wire [12:0]conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2;
    wire [12:0]conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2;
    wire [31:0]conv_core_inst_for_for_for_for_if_asn_6_itm_2;
    wire [31:0]conv_core_inst_for_for_for_for_if_asn_7_itm_2;
    wire nx63825z15, nx63825z14, nx63825z13, nx63825z12, nx63825z11, nx63825z10, 
         nx63825z9, nx63825z8, nx63825z7, nx63825z6, nx63825z5, nx63825z4, 
         nx63825z3, nx63825z2, nx63825z1;
    wire [31:31]conv_core_inst_z_out_4;
    wire \z_out_4(18)  , \z_out_4(19)  , \z_out_4(20)  , \z_out_4(21)  , 
         \z_out_4(22)  , \z_out_4(23)  , \z_out_4(24)  , \z_out_4(25)  , 
         \z_out_4(26)  , \z_out_4(27)  , \z_out_4(28)  , \z_out_4(29)  , 
         \z_out_4(30)  , \z_out_4(31)  , nx18281z15, nx18281z14, nx18281z13, 
         nx18281z12, nx18281z11, nx18281z10, nx18281z9, nx18281z8, nx18281z7, 
         nx18281z6, nx18281z5, nx18281z4, nx18281z3, nx18281z2, nx18281z1, 
         nx63825z63, nx63825z62, nx63825z61, nx63825z60, nx63825z59, nx63825z58, 
         nx63825z57, nx63825z56, nx63825z55, nx63825z54, nx63825z53, nx63825z52, 
         nx63825z51, nx63825z50, nx63825z49, nx63825z48, nx63825z47, nx63825z46, 
         nx63825z45, nx63825z44, nx63825z43, nx63825z42, nx63825z41, nx63825z40, 
         nx63825z39, nx63825z38, nx63825z37, nx63825z36, nx63825z35, nx63825z34, 
         nx63825z33, nx63825z32, nx63825z31, nx63825z30, nx63825z29, nx63825z28, 
         nx63825z27, nx63825z26, nx63825z25, nx63825z24, nx63825z23, nx63825z22, 
         nx63825z21, nx63825z20, nx63825z19, nx63825z18, nx63825z17, nx63825z16, 
         nx30685z34, nx30685z33, nx30685z32, nx30685z31, nx30685z30, nx30685z29, 
         nx30685z28, nx30685z27, nx30685z26, nx30685z25, nx30685z24, nx30685z23, 
         nx30685z22, nx30685z21, nx30685z20, nx30685z19, nx30685z18, nx30685z17, 
         nx30685z16, nx30685z15, nx30685z14, nx30685z13, nx30685z12, nx30685z11, 
         nx30685z10, nx30685z9, nx30685z8, nx30685z7, nx30685z6, nx30685z5, 
         nx30685z4, nx30685z3, nx30685z2, nx30685z1, nx18281z81, nx18281z80, 
         nx18281z79, nx18281z78, nx18281z77, nx18281z76, nx18281z75, nx18281z74, 
         nx18281z73, nx18281z72, nx18281z71, nx18281z70, nx18281z69, nx18281z68, 
         nx18281z67, nx18281z66, nx18281z65, nx18281z64, nx18281z63, nx18281z62, 
         nx18281z61, nx18281z60, nx18281z59, nx18281z58, nx18281z57, nx18281z56, 
         nx18281z55, nx18281z54, nx18281z53, nx18281z52, nx18281z51, nx18281z50, 
         nx18281z49, nx18281z48, nx18281z47, nx18281z46, nx18281z45, nx18281z44, 
         nx18281z43, nx18281z42, nx18281z41, nx18281z40, nx18281z39, nx18281z38, 
         nx18281z37, nx18281z36, nx18281z35, nx18281z34, \z_out_4(13)  , 
         \z_out_4(14)  , \z_out_4(15)  , \z_out_4(16)  , nx18281z33, nx18281z32, 
         nx18281z31, nx18281z30, nx18281z29, nx18281z28, nx18281z27, nx18281z26, 
         nx18281z25, nx18281z24, nx18281z23, nx18281z22, nx18281z21, nx18281z20, 
         nx18281z19, nx18281z18, nx18281z17, nx18281z16;
    wire \z_out_1(32)  ;
    wire nx49642z2, nx34566z1, nx49642z4, nx49641z2, nx49642z1, nx49641z3, 
         nx48653z2, nx49641z1, nx48653z3, nx48652z2, nx48653z1, nx48652z3, 
         nx48651z3, nx48652z1, nx48651z4, nx48650z2, nx48651z2, nx48650z3, 
         nx48649z2, nx48650z1, nx48649z3, nx48648z2, nx48649z1, nx48648z3, 
         nx48647z2, nx48648z1, nx48647z3, nx48646z2, nx48647z1, nx48646z3, 
         nx48645z2, nx48646z1, nx48645z3, nx48644z2, nx48645z1, nx48644z3, 
         nx47656z2, nx48644z1, nx47656z3, nx47655z2, nx47656z1, nx47655z3, 
         nx47654z3, nx47655z1, nx47654z4, nx47653z2, nx47654z2, nx47653z3, 
         nx47652z2, nx47653z1, nx47652z3, nx47651z2, nx47652z1, nx47651z3, 
         nx47650z2, nx47651z1, nx47650z3, nx47649z2, nx47650z1, nx47649z3, 
         nx47648z2, nx47649z1, nx47648z3, nx47647z2, nx47648z1, nx47647z3, 
         nx28341z2, nx47647z1, nx28341z3, nx28342z2, nx28341z1, nx28342z3, 
         nx28343z2, nx28342z1, nx28343z3, nx28344z2, nx28343z1, nx28344z3, 
         nx28345z2, nx28344z1, nx28345z3, nx28346z2, nx28345z1, nx28346z3, 
         nx28347z2, nx28346z1, nx28347z3, nx28348z2, nx28347z1, nx28348z3, 
         nx28349z2, nx28348z1, nx28349z3, nx28350z1, nx28349z1, nx28350z3, 
         not_fsm_output_5, nx50037z2, nx50037z1, nx50037z3, nx39519z4, nx39523z3, 
         nx39523z1, nx39523z2, nx39522z2, nx39518z4, nx39522z3, nx39521z3, 
         nx39521z2, nx39522z1, nx39520z3, nx39520z2, nx39521z1, nx39519z3, 
         nx39519z2, nx39520z1, nx39518z3, nx39518z2, nx39519z1, nx39517z5, 
         nx39517z2, nx39518z1, nx50045z2, nx39517z3, nx39517z1, nx48536z2, 
         nx60570z2, nx49524z2, nx48536z1, nx49525z2, nx49524z1, nx49526z2, 
         nx49525z1, nx49527z2, nx49526z1, nx49528z2, nx49527z1, nx49529z2, 
         nx49528z1, nx49530z2, nx49529z1, nx49531z2, nx49530z1, nx49532z2, 
         nx49531z1, nx49533z2, nx49532z1, nx50521z2, nx49533z1, nx50522z2, 
         nx50521z1, nx50523z2, nx50522z1, nx50524z2, nx50523z1, nx50525z2, 
         nx50524z1, nx50526z2, nx50525z1, nx50527z2, nx50526z1, nx50528z2, 
         nx50527z1, nx50529z2, nx50528z1, nx50530z2, nx50529z1, nx34270z2, 
         nx50530z1, nx34269z2, nx34270z1, nx34268z2, nx34269z1, nx34267z2, 
         nx34268z1, nx34266z2, nx34267z1, nx34265z2, nx34266z1, nx34264z2, 
         nx34265z1, nx34263z2, nx34264z1, nx34262z2, nx34263z1, nx34261z1, 
         nx34262z1, nx38873z2, nx38873z1, nx53949z2, nx53949z1, nx53948z2, 
         nx53948z1, nx34908z2, nx34908z1, nx34909z2, nx34909z1, nx34910z2, 
         nx34910z1, nx34911z2, nx34911z1, nx34912z2, nx34912z1, nx34913z2, 
         nx34913z1, nx34914z2, nx34914z1, nx34915z2, nx34915z1, nx34916z2, 
         nx34916z1, nx34917z1, nx7619z2;
    wire [31:0]conv_core_inst_for_for_for_for_acc_3_tmp;
    wire nx7619z1, nx7618z2, nx7618z1, nx6630z2, nx6630z1, nx6629z2, nx6629z1, 
         nx6628z2, nx6628z1, nx6627z2, nx6627z1, nx6626z2, nx6626z1, nx6625z2, 
         nx6625z1, nx6624z2, nx6624z1, nx6623z2, nx6623z1, nx6622z2, nx6622z1, 
         nx6621z2, nx6621z1, nx5633z2, nx5633z1, nx5632z2, nx5632z1, nx5631z2, 
         nx5631z1, nx5630z2, nx5630z1, nx5629z2, nx5629z1, nx5628z2, nx5628z1, 
         nx5627z2, nx5627z1, nx5626z2, nx5626z1, nx44834z2, nx44834z1, nx44835z2, 
         nx44835z1, nx8911z2, nx8911z1, nx8912z2, nx8912z1, nx8913z2, nx8913z1, 
         nx8914z2, nx8914z1, nx8915z2, nx8915z1, nx8916z2, 
         \for_for_for_acc_1_psp_sva_11n1s2(3)  , nx8916z1, nx8917z2, nx19541z2, 
         nx8917z1, nx8918z2, nx20538z2, nx8918z1, nx8919z2, nx12614z3, nx8919z1, 
         nx8920z1, nx64982z2;
    wire [31:0]conv_core_inst_jj_sva;
    wire \for_for_j_sva(30)  , nx64982z1, nx64981z2, \for_for_j_sva(29)  , 
         nx64981z1, nx63993z2, \for_for_j_sva(28)  , nx63993z1, nx63992z2, 
         \for_for_j_sva(27)  , nx63992z1, nx63991z2, \for_for_j_sva(26)  , 
         nx63991z1, nx63990z2, \for_for_j_sva(25)  , nx63990z1, nx63989z2, 
         \for_for_j_sva(24)  , nx63989z1, nx63988z2, \for_for_j_sva(23)  , 
         nx63988z1, nx63987z2, \for_for_j_sva(22)  , nx63987z1, nx63986z2, 
         \for_for_j_sva(21)  , nx63986z1, nx63985z2, \for_for_j_sva(20)  , 
         nx63985z1, nx63984z2, \for_for_j_sva(19)  , nx63984z1, nx62996z2, 
         \for_for_j_sva(18)  , nx62996z1, nx62995z2, \for_for_j_sva(17)  , 
         nx62995z1, nx62994z2, \for_for_j_sva(16)  , nx62994z1, nx62993z2, 
         \for_for_j_sva(15)  , nx62993z1, nx62992z2, \for_for_j_sva(14)  , 
         nx62992z1, nx62991z2, \for_for_j_sva(13)  , nx62991z1, nx62990z2, 
         \for_for_j_sva(12)  , nx62990z1, nx62989z2, \for_for_j_sva(11)  , 
         nx62989z1, nx62988z2, \for_for_j_sva(10)  , nx62988z1, nx62987z2, 
         \for_for_j_sva(9)  , nx62987z1, nx63175z2, \for_for_j_sva(8)  , 
         nx63175z1, nx63174z2, \for_for_j_sva(7)  , nx63174z1, nx63173z2, 
         \for_for_j_sva(6)  , nx63173z1, nx63172z2, \for_for_j_sva(5)  , 
         nx63172z1, nx63171z2, \for_for_j_sva(4)  , nx63171z1, nx63170z2, 
         \kernel_rsci_addr_d_0n0s2(3)  , nx63170z1, nx63169z2, 
         \for_for_for_for_n_4_0_sva(2)  , nx63169z1, nx63168z2, 
         \for_for_for_for_n_4_0_sva(1)  , nx63168z1, nx63167z2, 
         \for_for_for_for_n_4_0_sva(0)  , nx63167z1, nx63166z2, nx11961z2;
    wire [13:0]conv_core_inst_for_for_for_for_if_acc_psp_sva;
    wire \z_out_4(12)  , nx11961z1, nx11962z2, \z_out_4(11)  , nx11962z1, 
         nx11963z2, \z_out_4(10)  , nx11963z1, nx11964z2, \z_out_4(9)  , 
         nx11964z1, nx23668z2, \z_out_4(8)  , nx23668z1, nx23669z2, \z_out_4(7)  , 
         nx23669z1, nx23670z2, \z_out_4(6)  , nx23670z1, nx23671z2, \z_out_4(5)  , 
         nx23671z1, nx23672z2, \z_out_4(4)  , nx23672z1, nx23673z2, \z_out_4(3)  , 
         nx23673z1, nx23674z2, \z_out_4(2)  , nx23674z1, nx23675z2, \z_out_4(1)  , 
         nx23675z1, nx23676z2, \z_out_4(0)  , nx23676z1, nx23677z1, nx21390z2, 
         \z_out_2(0)  , \z_out_2(1)  , \z_out_2(2)  , \z_out_2(3)  , 
         \z_out_2(4)  , \z_out_2(5)  , \z_out_2(6)  , \z_out_2(7)  , 
         \z_out_2(8)  , \z_out_2(9)  , \z_out_2(10)  , \z_out_2(11)  , 
         \z_out_2(12)  , \z_out_2(13)  , \z_out_2(14)  , \z_out_2(15)  , 
         \z_out_2(16)  , \z_out_2(17)  , \z_out_2(18)  , \z_out_2(19)  , 
         \z_out_2(20)  , \z_out_2(21)  , \z_out_2(22)  , \z_out_2(23)  , 
         \z_out_2(24)  , \z_out_2(25)  , \z_out_2(26)  , \z_out_2(27)  , 
         \z_out_2(28)  , \z_out_2(29)  , \z_out_2(30)  ;
    wire [539:0] \$dummy ;




    inc_31_0 z_out_2_inc31_9 (.d ({\z_out_2(30)  ,\z_out_2(29)  ,\z_out_2(28)  ,
             \z_out_2(27)  ,\z_out_2(26)  ,\z_out_2(25)  ,\z_out_2(24)  ,
             \z_out_2(23)  ,\z_out_2(22)  ,\z_out_2(21)  ,\z_out_2(20)  ,
             \z_out_2(19)  ,\z_out_2(18)  ,\z_out_2(17)  ,\z_out_2(16)  ,
             \z_out_2(15)  ,\z_out_2(14)  ,\z_out_2(13)  ,\z_out_2(12)  ,
             \z_out_2(11)  ,\z_out_2(10)  ,\z_out_2(9)  ,\z_out_2(8)  ,
             \z_out_2(7)  ,\z_out_2(6)  ,\z_out_2(5)  ,\z_out_2(4)  ,
             \z_out_2(3)  ,\z_out_2(2)  ,\z_out_2(1)  ,\z_out_2(0)  }), .cout (
             nx21390z2), .\p_rows_rsc_z_int(30)   (p_nbus_rows_rsc_z_int[1]), .\p_fsm_output(9)   (
             \fsm_output(9)  ), .\p_fsm_output(0)   (\fsm_output(0)  ), .\p_for_i_sva(30)   (
             conv_core_inst_for_i_sva[26]), .px1533 (nx6185z1), .\p_rows_rsc_z_int(29)   (
             p_nbus_rows_rsc_z_int[2]), .\p_for_i_sva(29)   (
             conv_core_inst_for_i_sva[25]), .px1531 (nx6185z2), .\p_rows_rsc_z_int(28)   (
             p_nbus_rows_rsc_z_int[3]), .\p_for_i_sva(28)   (
             conv_core_inst_for_i_sva[24]), .px1529 (nx6185z3), .\p_rows_rsc_z_int(27)   (
             p_nbus_rows_rsc_z_int[4]), .\p_for_i_sva(27)   (
             conv_core_inst_for_i_sva[23]), .px1527 (nx6185z4), .\p_rows_rsc_z_int(26)   (
             p_nbus_rows_rsc_z_int[5]), .\p_for_i_sva(26)   (
             conv_core_inst_for_i_sva[22]), .px1525 (nx6185z5), .\p_rows_rsc_z_int(25)   (
             p_nbus_rows_rsc_z_int[6]), .\p_for_i_sva(25)   (
             conv_core_inst_for_i_sva[21]), .px1523 (nx6185z6), .\p_rows_rsc_z_int(24)   (
             p_nbus_rows_rsc_z_int[7]), .\p_for_i_sva(24)   (
             conv_core_inst_for_i_sva[20]), .px1521 (nx6185z7), .\p_rows_rsc_z_int(23)   (
             p_nbus_rows_rsc_z_int[8]), .\p_for_i_sva(23)   (
             conv_core_inst_for_i_sva[19]), .px1519 (nx6185z8), .\p_rows_rsc_z_int(22)   (
             p_nbus_rows_rsc_z_int[9]), .\p_for_i_sva(22)   (
             conv_core_inst_for_i_sva[18]), .px1517 (nx6185z9), .\p_rows_rsc_z_int(21)   (
             p_nbus_rows_rsc_z_int[10]), .\p_for_i_sva(21)   (
             conv_core_inst_for_i_sva[17]), .px1515 (nx6185z10), .\p_rows_rsc_z_int(20)   (
             p_nbus_rows_rsc_z_int[11]), .\p_for_i_sva(20)   (
             conv_core_inst_for_i_sva[16]), .px1513 (nx6185z11), .\p_rows_rsc_z_int(19)   (
             p_nbus_rows_rsc_z_int[12]), .\p_for_i_sva(19)   (
             conv_core_inst_for_i_sva[15]), .px1511 (nx6185z12), .\p_rows_rsc_z_int(18)   (
             p_nbus_rows_rsc_z_int[13]), .\p_for_i_sva(18)   (
             conv_core_inst_for_i_sva[14]), .px1509 (nx6185z13), .\p_rows_rsc_z_int(17)   (
             p_nbus_rows_rsc_z_int[14]), .\p_for_i_sva(17)   (
             conv_core_inst_for_i_sva[13]), .px1507 (nx6185z14), .\p_rows_rsc_z_int(16)   (
             p_nbus_rows_rsc_z_int[15]), .\p_for_i_sva(16)   (
             conv_core_inst_for_i_sva[12]), .px1505 (nx6185z15), .\p_rows_rsc_z_int(15)   (
             p_nbus_rows_rsc_z_int[16]), .\p_for_i_sva(15)   (
             conv_core_inst_for_i_sva[11]), .px1503 (nx6185z16), .\p_rows_rsc_z_int(14)   (
             p_nbus_rows_rsc_z_int[17]), .\p_for_i_sva(14)   (
             conv_core_inst_for_i_sva[10]), .px1501 (nx6185z17), .\p_rows_rsc_z_int(13)   (
             p_nbus_rows_rsc_z_int[18]), .\p_for_i_sva(13)   (
             conv_core_inst_for_i_sva[9]), .px1499 (nx6185z18), .\p_rows_rsc_z_int(12)   (
             p_nbus_rows_rsc_z_int[19]), .\p_for_i_sva(12)   (
             conv_core_inst_for_i_sva[8]), .px1497 (nx6185z19), .\p_rows_rsc_z_int(11)   (
             p_nbus_rows_rsc_z_int[20]), .\p_for_i_sva(11)   (
             conv_core_inst_for_i_sva[7]), .px1495 (nx6185z20), .\p_rows_rsc_z_int(10)   (
             p_nbus_rows_rsc_z_int[21]), .\p_for_i_sva(10)   (
             conv_core_inst_for_i_sva[6]), .px1493 (nx6185z21), .\p_rows_rsc_z_int(9)   (
             p_nbus_rows_rsc_z_int[22]), .\p_for_i_sva(9)   (
             conv_core_inst_for_i_sva[5]), .px1491 (nx6185z22), .\p_rows_rsc_z_int(8)   (
             p_nbus_rows_rsc_z_int[23]), .\p_for_i_sva(8)   (
             conv_core_inst_for_i_sva[4]), .px1489 (nx6185z23), .\p_rows_rsc_z_int(7)   (
             p_nbus_rows_rsc_z_int[24]), .\p_for_i_sva(7)   (
             conv_core_inst_for_i_sva[3]), .px1487 (nx6185z24), .\p_rows_rsc_z_int(6)   (
             p_nbus_rows_rsc_z_int[25]), .\p_for_i_sva(6)   (
             conv_core_inst_for_i_sva[2]), .px1485 (nx6185z25), .\p_rows_rsc_z_int(5)   (
             p_nbus_rows_rsc_z_int[26]), .\p_for_i_sva(5)   (
             conv_core_inst_for_i_sva[1]), .px1483 (nx6185z26), .\p_rows_rsc_z_int(4)   (
             p_nbus_rows_rsc_z_int[27]), .\p_for_i_sva(4)   (
             conv_core_inst_for_i_sva[0]), .px1481 (nx6185z27), .\p_rows_rsc_z_int(3)   (
             p_nbus_rows_rsc_z_int[28]), .\p_for_i_sva(3)   (
             conv_core_inst_for_i_sva[28]), .px1479 (nx6185z28), .\p_sortie_rsc_addr_1_0(2)   (
             \p_sortie_rsc_addr_1_0(2)  ), .\p_rows_rsc_z_int(2)   (
             p_nbus_rows_rsc_z_int[29]), .\p_fsm_output(8)   (\fsm_output(8)  )
             , .px1477 (nx6185z29), .\p_sortie_rsc_addr_1_0(1)   (
             \p_sortie_rsc_addr_1_0(1)  ), .\p_rows_rsc_z_int(1)   (
             p_nbus_rows_rsc_z_int[30]), .px1475 (nx6185z30), .\p_sortie_rsc_addr_1_0(0)   (
             \p_sortie_rsc_addr_1_0(0)  ), .\p_rows_rsc_z_int(0)   (
             p_nbus_rows_rsc_z_int[31]), .px1473 (nx6185z31)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_0 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[0]), .CI (px1140), .LI (
          nx23677z1)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_1 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[1]), .CI (nx23676z1), .LI (
          nx23676z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_2 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[2]), .CI (nx23675z1), .LI (
          nx23675z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_3 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[3]), .CI (nx23674z1), .LI (
          nx23674z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_4 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[4]), .CI (nx23673z1), .LI (
          nx23673z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_5 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[5]), .CI (nx23672z1), .LI (
          nx23672z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_6 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[6]), .CI (nx23671z1), .LI (
          nx23671z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_7 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[7]), .CI (nx23670z1), .LI (
          nx23670z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_8 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[8]), .CI (nx23669z1), .LI (
          nx23669z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_9 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[9]), .CI (nx23668z1), .LI (
          nx23668z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_10 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[10]), .CI (nx11964z1), .LI (
          nx11964z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_11 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[11]), .CI (nx11963z1), .LI (
          nx11963z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_12 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[12]), .CI (nx11962z1), .LI (
          nx11962z2)) ;
    XORCY for_for_for_for_if_acc_psp_sva_add14_0_xorcy_13 (.O (
          conv_core_inst_for_for_for_for_if_acc_psp_sva[13]), .CI (nx11961z1), .LI (
          nx11961z2)) ;
    XORCY jj_sva_add32_2_xorcy_0 (.O (conv_core_inst_jj_sva[0]), .CI (px1140), .LI (
          nx63166z2)) ;
    XORCY jj_sva_add32_2_xorcy_1 (.O (conv_core_inst_jj_sva[1]), .CI (nx63167z1)
          , .LI (nx63167z2)) ;
    XORCY jj_sva_add32_2_xorcy_2 (.O (conv_core_inst_jj_sva[2]), .CI (nx63168z1)
          , .LI (nx63168z2)) ;
    XORCY jj_sva_add32_2_xorcy_3 (.O (conv_core_inst_jj_sva[3]), .CI (nx63169z1)
          , .LI (nx63169z2)) ;
    XORCY jj_sva_add32_2_xorcy_4 (.O (conv_core_inst_jj_sva[4]), .CI (nx63170z1)
          , .LI (nx63170z2)) ;
    XORCY jj_sva_add32_2_xorcy_5 (.O (conv_core_inst_jj_sva[5]), .CI (nx63171z1)
          , .LI (nx63171z2)) ;
    XORCY jj_sva_add32_2_xorcy_6 (.O (conv_core_inst_jj_sva[6]), .CI (nx63172z1)
          , .LI (nx63172z2)) ;
    XORCY jj_sva_add32_2_xorcy_7 (.O (conv_core_inst_jj_sva[7]), .CI (nx63173z1)
          , .LI (nx63173z2)) ;
    XORCY jj_sva_add32_2_xorcy_8 (.O (conv_core_inst_jj_sva[8]), .CI (nx63174z1)
          , .LI (nx63174z2)) ;
    XORCY jj_sva_add32_2_xorcy_9 (.O (conv_core_inst_jj_sva[9]), .CI (nx63175z1)
          , .LI (nx63175z2)) ;
    XORCY jj_sva_add32_2_xorcy_10 (.O (conv_core_inst_jj_sva[10]), .CI (
          nx62987z1), .LI (nx62987z2)) ;
    XORCY jj_sva_add32_2_xorcy_11 (.O (conv_core_inst_jj_sva[11]), .CI (
          nx62988z1), .LI (nx62988z2)) ;
    XORCY jj_sva_add32_2_xorcy_12 (.O (conv_core_inst_jj_sva[12]), .CI (
          nx62989z1), .LI (nx62989z2)) ;
    XORCY jj_sva_add32_2_xorcy_13 (.O (conv_core_inst_jj_sva[13]), .CI (
          nx62990z1), .LI (nx62990z2)) ;
    XORCY jj_sva_add32_2_xorcy_14 (.O (conv_core_inst_jj_sva[14]), .CI (
          nx62991z1), .LI (nx62991z2)) ;
    XORCY jj_sva_add32_2_xorcy_15 (.O (conv_core_inst_jj_sva[15]), .CI (
          nx62992z1), .LI (nx62992z2)) ;
    XORCY jj_sva_add32_2_xorcy_16 (.O (conv_core_inst_jj_sva[16]), .CI (
          nx62993z1), .LI (nx62993z2)) ;
    XORCY jj_sva_add32_2_xorcy_17 (.O (conv_core_inst_jj_sva[17]), .CI (
          nx62994z1), .LI (nx62994z2)) ;
    XORCY jj_sva_add32_2_xorcy_18 (.O (conv_core_inst_jj_sva[18]), .CI (
          nx62995z1), .LI (nx62995z2)) ;
    XORCY jj_sva_add32_2_xorcy_19 (.O (conv_core_inst_jj_sva[19]), .CI (
          nx62996z1), .LI (nx62996z2)) ;
    XORCY jj_sva_add32_2_xorcy_20 (.O (conv_core_inst_jj_sva[20]), .CI (
          nx63984z1), .LI (nx63984z2)) ;
    XORCY jj_sva_add32_2_xorcy_21 (.O (conv_core_inst_jj_sva[21]), .CI (
          nx63985z1), .LI (nx63985z2)) ;
    XORCY jj_sva_add32_2_xorcy_22 (.O (conv_core_inst_jj_sva[22]), .CI (
          nx63986z1), .LI (nx63986z2)) ;
    XORCY jj_sva_add32_2_xorcy_23 (.O (conv_core_inst_jj_sva[23]), .CI (
          nx63987z1), .LI (nx63987z2)) ;
    XORCY jj_sva_add32_2_xorcy_24 (.O (conv_core_inst_jj_sva[24]), .CI (
          nx63988z1), .LI (nx63988z2)) ;
    XORCY jj_sva_add32_2_xorcy_25 (.O (conv_core_inst_jj_sva[25]), .CI (
          nx63989z1), .LI (nx63989z2)) ;
    XORCY jj_sva_add32_2_xorcy_26 (.O (conv_core_inst_jj_sva[26]), .CI (
          nx63990z1), .LI (nx63990z2)) ;
    XORCY jj_sva_add32_2_xorcy_27 (.O (conv_core_inst_jj_sva[27]), .CI (
          nx63991z1), .LI (nx63991z2)) ;
    XORCY jj_sva_add32_2_xorcy_28 (.O (conv_core_inst_jj_sva[28]), .CI (
          nx63992z1), .LI (nx63992z2)) ;
    XORCY jj_sva_add32_2_xorcy_29 (.O (conv_core_inst_jj_sva[29]), .CI (
          nx63993z1), .LI (nx63993z2)) ;
    XORCY jj_sva_add32_2_xorcy_30 (.O (conv_core_inst_jj_sva[30]), .CI (
          nx64981z1), .LI (nx64981z2)) ;
    XORCY jj_sva_add32_2_xorcy_31 (.O (conv_core_inst_jj_sva[31]), .CI (
          nx64982z1), .LI (nx64982z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_0 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[0]), .CI (px1140), .LI (
          nx8920z1)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_1 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[1]), .CI (nx8919z1), .LI (
          nx8919z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_2 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[2]), .CI (nx8918z1), .LI (
          nx8918z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_3 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[3]), .CI (nx8917z1), .LI (
          nx8917z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_4 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[4]), .CI (nx8916z1), .LI (
          nx8916z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_5 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[5]), .CI (nx8915z1), .LI (
          nx8915z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_6 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[6]), .CI (nx8914z1), .LI (
          nx8914z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_7 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[7]), .CI (nx8913z1), .LI (
          nx8913z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_8 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[8]), .CI (nx8912z1), .LI (
          nx8912z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_9 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[9]), .CI (nx8911z1), .LI (
          nx8911z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_10 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[10]), .CI (nx44835z1), .LI (
          nx44835z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_11 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[11]), .CI (nx44834z1), .LI (
          nx44834z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_12 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[12]), .CI (nx5626z1), .LI (
          nx5626z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_13 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[13]), .CI (nx5627z1), .LI (
          nx5627z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_14 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[14]), .CI (nx5628z1), .LI (
          nx5628z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_15 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[15]), .CI (nx5629z1), .LI (
          nx5629z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_16 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[16]), .CI (nx5630z1), .LI (
          nx5630z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_17 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[17]), .CI (nx5631z1), .LI (
          nx5631z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_18 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[18]), .CI (nx5632z1), .LI (
          nx5632z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_19 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[19]), .CI (nx5633z1), .LI (
          nx5633z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_20 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[20]), .CI (nx6621z1), .LI (
          nx6621z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_21 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[21]), .CI (nx6622z1), .LI (
          nx6622z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_22 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[22]), .CI (nx6623z1), .LI (
          nx6623z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_23 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[23]), .CI (nx6624z1), .LI (
          nx6624z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_24 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[24]), .CI (nx6625z1), .LI (
          nx6625z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_25 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[25]), .CI (nx6626z1), .LI (
          nx6626z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_26 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[26]), .CI (nx6627z1), .LI (
          nx6627z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_27 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[27]), .CI (nx6628z1), .LI (
          nx6628z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_28 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[28]), .CI (nx6629z1), .LI (
          nx6629z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_29 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[29]), .CI (nx6630z1), .LI (
          nx6630z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_30 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[30]), .CI (nx7618z1), .LI (
          nx7618z2)) ;
    XORCY for_for_for_for_acc_3_tmp_add32_3_xorcy_31 (.O (
          conv_core_inst_for_for_for_for_acc_3_tmp[31]), .CI (nx7619z1), .LI (
          nx7619z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_0 (.O (p_nbus_image_rsc_addr_1_0[0]), 
          .CI (px1140), .LI (nx34917z1)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_1 (.O (p_nbus_image_rsc_addr_1_0[1]), 
          .CI (nx34916z1), .LI (nx34916z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_2 (.O (p_nbus_image_rsc_addr_1_0[2]), 
          .CI (nx34915z1), .LI (nx34915z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_3 (.O (p_nbus_image_rsc_addr_1_0[3]), 
          .CI (nx34914z1), .LI (nx34914z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_4 (.O (p_nbus_image_rsc_addr_1_0[4]), 
          .CI (nx34913z1), .LI (nx34913z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_5 (.O (p_nbus_image_rsc_addr_1_0[5]), 
          .CI (nx34912z1), .LI (nx34912z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_6 (.O (p_nbus_image_rsc_addr_1_0[6]), 
          .CI (nx34911z1), .LI (nx34911z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_7 (.O (p_nbus_image_rsc_addr_1_0[7]), 
          .CI (nx34910z1), .LI (nx34910z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_8 (.O (p_nbus_image_rsc_addr_1_0[8]), 
          .CI (nx34909z1), .LI (nx34909z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_9 (.O (p_nbus_image_rsc_addr_1_0[9]), 
          .CI (nx34908z1), .LI (nx34908z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_10 (.O (p_nbus_image_rsc_addr_1_0[10])
          , .CI (nx53948z1), .LI (nx53948z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_11 (.O (p_nbus_image_rsc_addr_1_0[11])
          , .CI (nx53949z1), .LI (nx53949z2)) ;
    XORCY image_rsci_addr_d_add13_4_xorcy_12 (.O (p_nbus_image_rsc_addr_1_0[12])
          , .CI (nx38873z1), .LI (nx38873z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_30 (.O (nx60570z2), .CI (
          nx48536z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[30]), .S (
          nx48536z2)) ;
    GND ps_gnd (.G (nx39517z1)) ;
    VCC ps_vcc (.P (nx39517z3)) ;
    XORCY xorcy_0_0 (.O (p_nbus_kernel_rsc_addr_1_0[0]), .CI (nx39517z1), .LI (
          nx50045z2)) ;
    XORCY xorcy_0_1 (.O (p_nbus_kernel_rsc_addr_1_0[1]), .CI (nx39517z1), .LI (
          nx39517z5)) ;
    XORCY xorcy_0_2 (.O (p_nbus_kernel_rsc_addr_1_0[2]), .CI (nx39518z1), .LI (
          nx39518z3)) ;
    XORCY xorcy_0_3 (.O (p_nbus_kernel_rsc_addr_1_0[3]), .CI (nx39519z1), .LI (
          nx39519z3)) ;
    XORCY xorcy_0_4 (.O (p_nbus_kernel_rsc_addr_1_0[4]), .CI (nx39520z1), .LI (
          nx39520z3)) ;
    XORCY xorcy_0_5 (.O (p_nbus_kernel_rsc_addr_1_0[5]), .CI (nx39521z1), .LI (
          nx39521z3)) ;
    (* HLUTNM = "conv_core_inst_modgen_adderblock_slut_0_6" *)
    LUT4 slut_0_6 (.O (nx39522z3), .I0 (nx39518z4), .I1 (nx39517z1), .I2 (
         nx39517z3), .I3 (nx39522z2)) ;
         defparam slut_0_6.INIT = 16'h6996;
    (* HLUTNM = "conv_core_inst_modgen_adderblock_slut_0_6" *)
    LUT3 clut_0_6 (.O (nx39523z2), .I0 (nx39518z4), .I1 (nx39517z1), .I2 (
         nx39517z3)) ;
         defparam clut_0_6.INIT = 8'hE8;
    XORCY xorcy_0_6 (.O (p_nbus_kernel_rsc_addr_1_0[6]), .CI (nx39522z1), .LI (
          nx39522z3)) ;
    (* HLUTNM = "conv_core_inst_modgen_adderblock_slut_0_7" *)
    LUT4 slut_0_7 (.O (nx39523z3), .I0 (nx39519z4), .I1 (nx39517z1), .I2 (
         nx39517z3), .I3 (nx39523z2)) ;
         defparam slut_0_7.INIT = 16'h6996;
    (* HLUTNM = "conv_core_inst_modgen_adderblock_slut_0_7" *)
    LUT3 clut_0_7 (.O (nx50037z3), .I0 (nx39519z4), .I1 (nx39517z1), .I2 (
         nx39517z3)) ;
         defparam clut_0_7.INIT = 8'hE8;
    XORCY xorcy_0_7 (.O (p_nbus_kernel_rsc_addr_1_0[7]), .CI (nx39523z1), .LI (
          nx39523z3)) ;
    XORCY xorcy_0_8 (.O (p_nbus_kernel_rsc_addr_1_0[8]), .CI (nx50037z1), .LI (
          nx50037z2)) ;
    XORCY z_out_1_add34_7_xorcy_0 (.O (p_nbus_sortie_rsc_data_in_1_0[0]), .CI (
          not_fsm_output_5), .LI (nx28350z3)) ;
    XORCY z_out_1_add34_7_xorcy_1 (.O (p_nbus_sortie_rsc_data_in_1_0[1]), .CI (
          nx28349z1), .LI (nx28349z3)) ;
    XORCY z_out_1_add34_7_xorcy_2 (.O (p_nbus_sortie_rsc_data_in_1_0[2]), .CI (
          nx28348z1), .LI (nx28348z3)) ;
    XORCY z_out_1_add34_7_xorcy_3 (.O (p_nbus_sortie_rsc_data_in_1_0[3]), .CI (
          nx28347z1), .LI (nx28347z3)) ;
    XORCY z_out_1_add34_7_xorcy_4 (.O (p_nbus_sortie_rsc_data_in_1_0[4]), .CI (
          nx28346z1), .LI (nx28346z3)) ;
    XORCY z_out_1_add34_7_xorcy_5 (.O (p_nbus_sortie_rsc_data_in_1_0[5]), .CI (
          nx28345z1), .LI (nx28345z3)) ;
    XORCY z_out_1_add34_7_xorcy_6 (.O (p_nbus_sortie_rsc_data_in_1_0[6]), .CI (
          nx28344z1), .LI (nx28344z3)) ;
    XORCY z_out_1_add34_7_xorcy_7 (.O (p_nbus_sortie_rsc_data_in_1_0[7]), .CI (
          nx28343z1), .LI (nx28343z3)) ;
    XORCY z_out_1_add34_7_xorcy_8 (.O (p_nbus_sortie_rsc_data_in_1_0[8]), .CI (
          nx28342z1), .LI (nx28342z3)) ;
    XORCY z_out_1_add34_7_xorcy_9 (.O (p_nbus_sortie_rsc_data_in_1_0[9]), .CI (
          nx28341z1), .LI (nx28341z3)) ;
    XORCY z_out_1_add34_7_xorcy_10 (.O (p_nbus_sortie_rsc_data_in_1_0[10]), .CI (
          nx47647z1), .LI (nx47647z3)) ;
    XORCY z_out_1_add34_7_xorcy_11 (.O (p_nbus_sortie_rsc_data_in_1_0[11]), .CI (
          nx47648z1), .LI (nx47648z3)) ;
    XORCY z_out_1_add34_7_xorcy_12 (.O (p_nbus_sortie_rsc_data_in_1_0[12]), .CI (
          nx47649z1), .LI (nx47649z3)) ;
    XORCY z_out_1_add34_7_xorcy_13 (.O (p_nbus_sortie_rsc_data_in_1_0[13]), .CI (
          nx47650z1), .LI (nx47650z3)) ;
    XORCY z_out_1_add34_7_xorcy_14 (.O (p_nbus_sortie_rsc_data_in_1_0[14]), .CI (
          nx47651z1), .LI (nx47651z3)) ;
    XORCY z_out_1_add34_7_xorcy_15 (.O (p_nbus_sortie_rsc_data_in_1_0[15]), .CI (
          nx47652z1), .LI (nx47652z3)) ;
    XORCY z_out_1_add34_7_xorcy_16 (.O (p_nbus_sortie_rsc_data_in_1_0[16]), .CI (
          nx47653z1), .LI (nx47653z3)) ;
    XORCY z_out_1_add34_7_xorcy_17 (.O (p_nbus_sortie_rsc_data_in_1_0[17]), .CI (
          nx47654z2), .LI (nx47654z4)) ;
    XORCY z_out_1_add34_7_xorcy_18 (.O (p_nbus_sortie_rsc_data_in_1_0[18]), .CI (
          nx47655z1), .LI (nx47655z3)) ;
    XORCY z_out_1_add34_7_xorcy_19 (.O (p_nbus_sortie_rsc_data_in_1_0[19]), .CI (
          nx47656z1), .LI (nx47656z3)) ;
    XORCY z_out_1_add34_7_xorcy_20 (.O (p_nbus_sortie_rsc_data_in_1_0[20]), .CI (
          nx48644z1), .LI (nx48644z3)) ;
    XORCY z_out_1_add34_7_xorcy_21 (.O (p_nbus_sortie_rsc_data_in_1_0[21]), .CI (
          nx48645z1), .LI (nx48645z3)) ;
    XORCY z_out_1_add34_7_xorcy_22 (.O (p_nbus_sortie_rsc_data_in_1_0[22]), .CI (
          nx48646z1), .LI (nx48646z3)) ;
    XORCY z_out_1_add34_7_xorcy_23 (.O (p_nbus_sortie_rsc_data_in_1_0[23]), .CI (
          nx48647z1), .LI (nx48647z3)) ;
    XORCY z_out_1_add34_7_xorcy_24 (.O (p_nbus_sortie_rsc_data_in_1_0[24]), .CI (
          nx48648z1), .LI (nx48648z3)) ;
    XORCY z_out_1_add34_7_xorcy_25 (.O (p_nbus_sortie_rsc_data_in_1_0[25]), .CI (
          nx48649z1), .LI (nx48649z3)) ;
    XORCY z_out_1_add34_7_xorcy_26 (.O (p_nbus_sortie_rsc_data_in_1_0[26]), .CI (
          nx48650z1), .LI (nx48650z3)) ;
    XORCY z_out_1_add34_7_xorcy_27 (.O (p_nbus_sortie_rsc_data_in_1_0[27]), .CI (
          nx48651z2), .LI (nx48651z4)) ;
    XORCY z_out_1_add34_7_xorcy_28 (.O (p_nbus_sortie_rsc_data_in_1_0[28]), .CI (
          nx48652z1), .LI (nx48652z3)) ;
    XORCY z_out_1_add34_7_xorcy_29 (.O (p_nbus_sortie_rsc_data_in_1_0[29]), .CI (
          nx48653z1), .LI (nx48653z3)) ;
    XORCY z_out_1_add34_7_xorcy_30 (.O (p_nbus_sortie_rsc_data_in_1_0[30]), .CI (
          nx49641z1), .LI (nx49641z3)) ;
    XORCY z_out_1_add34_7_xorcy_31 (.O (p_nbus_sortie_rsc_data_in_1_0[31]), .CI (
          nx49642z1), .LI (nx49642z4)) ;
    XORCY z_out_1_add34_7_xorcy_32 (.O (\z_out_1(32)  ), .CI (nx34566z1), .LI (
          nx49642z4)) ;
    FDRE \reg_rows_1_sva_2(31)  (.Q (conv_core_inst_rows_1_sva_2[0]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[0]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(30)  (.Q (conv_core_inst_rows_1_sva_2[1]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[1]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(29)  (.Q (conv_core_inst_rows_1_sva_2[2]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[2]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(28)  (.Q (conv_core_inst_rows_1_sva_2[3]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[3]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(27)  (.Q (conv_core_inst_rows_1_sva_2[4]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[4]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(26)  (.Q (conv_core_inst_rows_1_sva_2[5]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[5]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(25)  (.Q (conv_core_inst_rows_1_sva_2[6]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[6]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(24)  (.Q (conv_core_inst_rows_1_sva_2[7]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[7]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(23)  (.Q (conv_core_inst_rows_1_sva_2[8]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[8]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(22)  (.Q (conv_core_inst_rows_1_sva_2[9]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[9]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(21)  (.Q (conv_core_inst_rows_1_sva_2[10]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[10]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(20)  (.Q (conv_core_inst_rows_1_sva_2[11]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[11]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(19)  (.Q (conv_core_inst_rows_1_sva_2[12]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[12]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(18)  (.Q (conv_core_inst_rows_1_sva_2[13]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[13]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(17)  (.Q (conv_core_inst_rows_1_sva_2[14]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[14]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(16)  (.Q (conv_core_inst_rows_1_sva_2[15]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[15]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(15)  (.Q (conv_core_inst_rows_1_sva_2[16]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[16]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(14)  (.Q (conv_core_inst_rows_1_sva_2[17]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[17]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(13)  (.Q (conv_core_inst_rows_1_sva_2[18]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[18]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(12)  (.Q (conv_core_inst_rows_1_sva_2[19]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[19]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(11)  (.Q (conv_core_inst_rows_1_sva_2[20]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[20]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(10)  (.Q (conv_core_inst_rows_1_sva_2[21]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[21]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(9)  (.Q (conv_core_inst_rows_1_sva_2[22]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[22]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(8)  (.Q (conv_core_inst_rows_1_sva_2[23]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[23]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(7)  (.Q (conv_core_inst_rows_1_sva_2[24]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[24]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(6)  (.Q (conv_core_inst_rows_1_sva_2[25]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[25]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(5)  (.Q (conv_core_inst_rows_1_sva_2[26]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[26]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(4)  (.Q (conv_core_inst_rows_1_sva_2[27]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[27]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(3)  (.Q (conv_core_inst_rows_1_sva_2[28]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[28]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(2)  (.Q (conv_core_inst_rows_1_sva_2[29]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[29]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(1)  (.Q (conv_core_inst_rows_1_sva_2[30]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[30]), .R (
         p_rst_int)) ;
    FDRE \reg_rows_1_sva_2(0)  (.Q (conv_core_inst_rows_1_sva_2[31]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_rows_rsc_z_int[31]), .R (
         p_rst_int)) ;
    FDRE \reg_for_i_sva(31)  (.Q (conv_core_inst_for_i_sva[27]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx65146z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(30)  (.Q (conv_core_inst_for_i_sva[26]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx64149z2), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(29)  (.Q (conv_core_inst_for_i_sva[25]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx62153z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(28)  (.Q (conv_core_inst_for_i_sva[24]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx61156z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(27)  (.Q (conv_core_inst_for_i_sva[23]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx60159z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(26)  (.Q (conv_core_inst_for_i_sva[22]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx59162z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(25)  (.Q (conv_core_inst_for_i_sva[21]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx58165z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(24)  (.Q (conv_core_inst_for_i_sva[20]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx57168z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(23)  (.Q (conv_core_inst_for_i_sva[19]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx56171z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(22)  (.Q (conv_core_inst_for_i_sva[18]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx55174z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(21)  (.Q (conv_core_inst_for_i_sva[17]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx54177z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(20)  (.Q (conv_core_inst_for_i_sva[16]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx53180z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(19)  (.Q (conv_core_inst_for_i_sva[15]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx51184z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(18)  (.Q (conv_core_inst_for_i_sva[14]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx50187z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(17)  (.Q (conv_core_inst_for_i_sva[13]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx49190z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(16)  (.Q (conv_core_inst_for_i_sva[12]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx48193z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(15)  (.Q (conv_core_inst_for_i_sva[11]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx47196z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(14)  (.Q (conv_core_inst_for_i_sva[10]), .C (p_clk_int)
         , .CE (nx64149z1), .D (nx46199z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(13)  (.Q (conv_core_inst_for_i_sva[9]), .C (p_clk_int), 
         .CE (nx64149z1), .D (nx45202z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(12)  (.Q (conv_core_inst_for_i_sva[8]), .C (p_clk_int), 
         .CE (nx64149z1), .D (nx44205z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(11)  (.Q (conv_core_inst_for_i_sva[7]), .C (p_clk_int), 
         .CE (nx64149z1), .D (nx43208z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(10)  (.Q (conv_core_inst_for_i_sva[6]), .C (p_clk_int), 
         .CE (nx64149z1), .D (nx42211z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(9)  (.Q (conv_core_inst_for_i_sva[5]), .C (p_clk_int), .CE (
         nx64149z1), .D (nx42669z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(8)  (.Q (conv_core_inst_for_i_sva[4]), .C (p_clk_int), .CE (
         nx64149z1), .D (nx43666z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(7)  (.Q (conv_core_inst_for_i_sva[3]), .C (p_clk_int), .CE (
         nx64149z1), .D (nx44663z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(6)  (.Q (conv_core_inst_for_i_sva[2]), .C (p_clk_int), .CE (
         nx64149z1), .D (nx45660z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(5)  (.Q (conv_core_inst_for_i_sva[1]), .C (p_clk_int), .CE (
         nx64149z1), .D (nx46657z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(4)  (.Q (conv_core_inst_for_i_sva[0]), .C (p_clk_int), .CE (
         nx64149z1), .D (nx47654z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(3)  (.Q (conv_core_inst_for_i_sva[28]), .C (p_clk_int), 
         .CE (nx64149z1), .D (nx48651z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(2)  (.Q (conv_core_inst_for_i_sva[29]), .C (p_clk_int), 
         .CE (nx64149z1), .D (nx49648z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(1)  (.Q (conv_core_inst_for_i_sva[30]), .C (p_clk_int), 
         .CE (nx64149z1), .D (nx50645z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_sva(0)  (.Q (conv_core_inst_for_i_sva[31]), .C (p_clk_int), 
         .CE (nx64149z1), .D (nx51642z1), .R (p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(31)  (.Q (conv_core_inst_cols_1_sva_1[0]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[0]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(30)  (.Q (conv_core_inst_cols_1_sva_1[1]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[1]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(29)  (.Q (conv_core_inst_cols_1_sva_1[2]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[2]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(28)  (.Q (conv_core_inst_cols_1_sva_1[3]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[3]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(27)  (.Q (conv_core_inst_cols_1_sva_1[4]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[4]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(26)  (.Q (conv_core_inst_cols_1_sva_1[5]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[5]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(25)  (.Q (conv_core_inst_cols_1_sva_1[6]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[6]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(24)  (.Q (conv_core_inst_cols_1_sva_1[7]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[7]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(23)  (.Q (conv_core_inst_cols_1_sva_1[8]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[8]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(22)  (.Q (conv_core_inst_cols_1_sva_1[9]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[9]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(21)  (.Q (conv_core_inst_cols_1_sva_1[10]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[10]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(20)  (.Q (conv_core_inst_cols_1_sva_1[11]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[11]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(19)  (.Q (conv_core_inst_cols_1_sva_1[12]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[12]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(18)  (.Q (conv_core_inst_cols_1_sva_1[13]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[13]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(17)  (.Q (conv_core_inst_cols_1_sva_1[14]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[14]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(16)  (.Q (conv_core_inst_cols_1_sva_1[15]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[15]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(15)  (.Q (conv_core_inst_cols_1_sva_1[16]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[16]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(14)  (.Q (conv_core_inst_cols_1_sva_1[17]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[17]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(13)  (.Q (conv_core_inst_cols_1_sva_1[18]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[18]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(12)  (.Q (conv_core_inst_cols_1_sva_1[19]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[19]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(11)  (.Q (conv_core_inst_cols_1_sva_1[20]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[20]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(10)  (.Q (conv_core_inst_cols_1_sva_1[21]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[21]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(9)  (.Q (conv_core_inst_cols_1_sva_1[22]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[22]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(8)  (.Q (conv_core_inst_cols_1_sva_1[23]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[23]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(7)  (.Q (conv_core_inst_cols_1_sva_1[24]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[24]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(6)  (.Q (conv_core_inst_cols_1_sva_1[25]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[25]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(5)  (.Q (conv_core_inst_cols_1_sva_1[26]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[26]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(4)  (.Q (conv_core_inst_cols_1_sva_1[27]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[27]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(3)  (.Q (conv_core_inst_cols_1_sva_1[28]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[28]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(2)  (.Q (conv_core_inst_cols_1_sva_1[29]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[29]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(1)  (.Q (conv_core_inst_cols_1_sva_1[30]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[30]), .R (
         p_rst_int)) ;
    FDRE \reg_cols_1_sva_1(0)  (.Q (conv_core_inst_cols_1_sva_1[31]), .C (
         p_clk_int), .CE (nx9631z1), .D (p_nbus_cols_rsc_z_int[31]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_j_sva(31)  (.Q (\for_for_j_sva(31)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx53153z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(30)  (.Q (\for_for_j_sva(30)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx52156z2), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(29)  (.Q (\for_for_j_sva(29)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx50160z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(28)  (.Q (\for_for_j_sva(28)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx49163z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(27)  (.Q (\for_for_j_sva(27)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx48166z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(26)  (.Q (\for_for_j_sva(26)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx47169z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(25)  (.Q (\for_for_j_sva(25)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx46172z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(24)  (.Q (\for_for_j_sva(24)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx45175z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(23)  (.Q (\for_for_j_sva(23)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx44178z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(22)  (.Q (\for_for_j_sva(22)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx43181z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(21)  (.Q (\for_for_j_sva(21)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx42184z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(20)  (.Q (\for_for_j_sva(20)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx41187z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(19)  (.Q (\for_for_j_sva(19)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx39191z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(18)  (.Q (\for_for_j_sva(18)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx38194z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(17)  (.Q (\for_for_j_sva(17)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx37197z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(16)  (.Q (\for_for_j_sva(16)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx36200z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(15)  (.Q (\for_for_j_sva(15)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx35203z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(14)  (.Q (\for_for_j_sva(14)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx34206z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(13)  (.Q (\for_for_j_sva(13)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx33209z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(12)  (.Q (\for_for_j_sva(12)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx32212z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(11)  (.Q (\for_for_j_sva(11)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx31215z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(10)  (.Q (\for_for_j_sva(10)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx30218z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(9)  (.Q (\for_for_j_sva(9)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx24210z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(8)  (.Q (\for_for_j_sva(8)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx25207z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(7)  (.Q (\for_for_j_sva(7)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx26204z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(6)  (.Q (\for_for_j_sva(6)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx27201z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(5)  (.Q (\for_for_j_sva(5)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx28198z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(4)  (.Q (\for_for_j_sva(4)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx29195z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(3)  (.Q (\for_for_j_sva(3)  ), .C (p_clk_int), .CE (
         nx52156z1), .D (nx30192z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(2)  (.Q (\p_sortie_rsc_addr_1_0(2)  ), .C (p_clk_int
         ), .CE (nx52156z1), .D (nx31189z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(1)  (.Q (\p_sortie_rsc_addr_1_0(1)  ), .C (p_clk_int
         ), .CE (nx52156z1), .D (nx32186z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_sva(0)  (.Q (\p_sortie_rsc_addr_1_0(0)  ), .C (p_clk_int
         ), .CE (nx52156z1), .D (nx33183z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(13)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[0]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[13]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(12)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[1]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[12]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(11)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[2]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[11]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(10)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[3]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[10]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(9)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[4]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[9]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(8)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[5]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[8]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(7)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[6]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[7]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(6)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[7]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[6]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(5)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[8]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[5]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(4)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[9]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[4]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(3)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[10]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[3]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(2)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[11]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[2]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(1)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[12]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[1]
         ), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_acc_psp_sva_1(0)  (.Q (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[13]), .C (p_clk_int), .CE (
         not_fsm_output_4), .D (conv_core_inst_for_for_for_for_if_acc_psp_sva[0]
         ), .R (p_rst_int)) ;
    FDRE reg_for_for_for_for_slc_for_for_for_for_acc_5_itm (.Q (
         for_for_for_for_slc_for_for_for_for_acc_5_itm), .C (p_clk_int), .CE (
         \fsm_output(3)  ), .D (nx12614z1), .R (p_rst_int)) ;
    FDRE reg_for_for_for_for_if_for_for_for_for_if_and_2_itm (.Q (
         for_for_for_for_if_for_for_for_for_if_and_2_itm), .C (p_clk_int), .CE (
         \fsm_output(3)  ), .D (nx60570z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva_3(4)  (.Q (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[0]), .C (p_clk_int), .CE (
         \fsm_output(3)  ), .D (nx20393z2), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva_3(3)  (.Q (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[1]), .C (p_clk_int), .CE (
         \fsm_output(3)  ), .D (nx18544z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva_3(2)  (.Q (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[2]), .C (p_clk_int), .CE (
         \fsm_output(3)  ), .D (nx19541z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva_3(1)  (.Q (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[3]), .C (p_clk_int), .CE (
         \fsm_output(3)  ), .D (nx20538z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva_3(0)  (.Q (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[4]), .C (p_clk_int), .CE (
         \fsm_output(3)  ), .D (nx12614z2), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_m_4_0_sva_4(4)  (.Q (nx20393z3), .C (p_clk_int), .CE (
         nx21003z1), .D (nx24991z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_m_4_0_sva_4(3)  (.Q (nx18544z2), .C (p_clk_int), .CE (
         nx21003z1), .D (nx23994z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_m_4_0_sva_4(2)  (.Q (nx19541z2), .C (p_clk_int), .CE (
         nx21003z1), .D (nx22997z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_m_4_0_sva_4(1)  (.Q (nx20538z2), .C (p_clk_int), .CE (
         nx21003z1), .D (nx22000z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_m_4_0_sva_4(0)  (.Q (nx12614z3), .C (p_clk_int), .CE (
         nx21003z1), .D (nx21003z2), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_acc_1_psp_sva(4)  (.Q (nx39520z4), .C (p_clk_int), .CE (
         nx59318z1), .D (nx55330z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_acc_1_psp_sva(3)  (.Q (nx39519z4), .C (p_clk_int), .CE (
         nx59318z1), .D (nx56327z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_acc_1_psp_sva(2)  (.Q (nx39518z4), .C (p_clk_int), .CE (
         nx59318z1), .D (nx57324z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_acc_1_psp_sva(1)  (.Q (nx39517z6), .C (p_clk_int), .CE (
         nx59318z1), .D (nx58321z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_acc_1_psp_sva(0)  (.Q (nx39517z4), .C (p_clk_int), .CE (
         nx59318z1), .D (nx12614z3), .R (p_rst_int)) ;
    LUT4 ix39521z28345 (.O (nx39521z3), .I0 (nx39517z6), .I1 (nx39520z4), .I2 (
         nx39517z3), .I3 (nx39521z2)) ;
         defparam ix39521z28345.INIT = 16'h6996;
    LUT3 ix39522z1546 (.O (nx39522z2), .I0 (nx39517z6), .I1 (nx39520z4), .I2 (
         nx39517z3)) ;
         defparam ix39522z1546.INIT = 8'hE8;
    LUT4 ix50037z28344 (.O (nx50037z2), .I0 (nx39520z4), .I1 (nx39517z1), .I2 (
         nx39517z3), .I3 (nx50037z3)) ;
         defparam ix50037z28344.INIT = 16'h6996;
    LUT2 ix23677z1320 (.O (nx23677z1), .I0 (\z_out_4(0)  ), .I1 (
         \for_for_j_sva(3)  )) ;
         defparam ix23677z1320.INIT = 4'h6;
    LUT2 ix23676z1320 (.O (nx23676z2), .I0 (\z_out_4(1)  ), .I1 (
         \for_for_j_sva(4)  )) ;
         defparam ix23676z1320.INIT = 4'h6;
    LUT2 ix23675z1320 (.O (nx23675z2), .I0 (\z_out_4(2)  ), .I1 (
         \for_for_j_sva(5)  )) ;
         defparam ix23675z1320.INIT = 4'h6;
    LUT2 ix23674z1320 (.O (nx23674z2), .I0 (\z_out_4(3)  ), .I1 (
         \for_for_j_sva(6)  )) ;
         defparam ix23674z1320.INIT = 4'h6;
    LUT2 ix23673z1320 (.O (nx23673z2), .I0 (\z_out_4(4)  ), .I1 (
         \for_for_j_sva(7)  )) ;
         defparam ix23673z1320.INIT = 4'h6;
    LUT2 ix23672z1320 (.O (nx23672z2), .I0 (\z_out_4(5)  ), .I1 (
         \for_for_j_sva(8)  )) ;
         defparam ix23672z1320.INIT = 4'h6;
    LUT2 ix23671z1320 (.O (nx23671z2), .I0 (\z_out_4(6)  ), .I1 (
         \for_for_j_sva(9)  )) ;
         defparam ix23671z1320.INIT = 4'h6;
    LUT2 ix23670z1320 (.O (nx23670z2), .I0 (\z_out_4(7)  ), .I1 (
         \for_for_j_sva(10)  )) ;
         defparam ix23670z1320.INIT = 4'h6;
    LUT2 ix23669z1320 (.O (nx23669z2), .I0 (\z_out_4(8)  ), .I1 (
         \for_for_j_sva(11)  )) ;
         defparam ix23669z1320.INIT = 4'h6;
    LUT2 ix23668z1320 (.O (nx23668z2), .I0 (\z_out_4(9)  ), .I1 (
         \for_for_j_sva(12)  )) ;
         defparam ix23668z1320.INIT = 4'h6;
    LUT2 ix11964z1320 (.O (nx11964z2), .I0 (\z_out_4(10)  ), .I1 (
         \for_for_j_sva(13)  )) ;
         defparam ix11964z1320.INIT = 4'h6;
    LUT2 ix11963z1320 (.O (nx11963z2), .I0 (\z_out_4(11)  ), .I1 (
         \for_for_j_sva(14)  )) ;
         defparam ix11963z1320.INIT = 4'h6;
    LUT2 ix11962z1320 (.O (nx11962z2), .I0 (\z_out_4(12)  ), .I1 (
         \for_for_j_sva(15)  )) ;
         defparam ix11962z1320.INIT = 4'h6;
    LUT2 ix11961z1320 (.O (nx11961z2), .I0 (\z_out_4(13)  ), .I1 (
         \for_for_j_sva(16)  )) ;
         defparam ix11961z1320.INIT = 4'h6;
    LUT2 ix63166z1320 (.O (nx63166z2), .I0 (\for_for_for_for_n_4_0_sva(0)  ), .I1 (
         \p_sortie_rsc_addr_1_0(0)  )) ;
         defparam ix63166z1320.INIT = 4'h6;
    LUT2 ix63167z1320 (.O (nx63167z2), .I0 (\for_for_for_for_n_4_0_sva(1)  ), .I1 (
         \p_sortie_rsc_addr_1_0(1)  )) ;
         defparam ix63167z1320.INIT = 4'h6;
    LUT2 ix63168z1320 (.O (nx63168z2), .I0 (\for_for_for_for_n_4_0_sva(2)  ), .I1 (
         \p_sortie_rsc_addr_1_0(2)  )) ;
         defparam ix63168z1320.INIT = 4'h6;
    LUT3 ix63170z1419 (.O (nx63170z2), .I0 (\for_for_j_sva(4)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63170z1419.INIT = 8'h69;
    LUT3 ix63171z1419 (.O (nx63171z2), .I0 (\for_for_j_sva(5)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63171z1419.INIT = 8'h69;
    LUT3 ix63172z1419 (.O (nx63172z2), .I0 (\for_for_j_sva(6)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63172z1419.INIT = 8'h69;
    LUT3 ix63173z1419 (.O (nx63173z2), .I0 (\for_for_j_sva(7)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63173z1419.INIT = 8'h69;
    LUT3 ix63174z1419 (.O (nx63174z2), .I0 (\for_for_j_sva(8)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63174z1419.INIT = 8'h69;
    LUT3 ix63175z1419 (.O (nx63175z2), .I0 (\for_for_j_sva(9)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63175z1419.INIT = 8'h69;
    LUT3 ix62987z1419 (.O (nx62987z2), .I0 (\for_for_j_sva(10)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62987z1419.INIT = 8'h69;
    LUT3 ix62988z1419 (.O (nx62988z2), .I0 (\for_for_j_sva(11)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62988z1419.INIT = 8'h69;
    LUT3 ix62989z1419 (.O (nx62989z2), .I0 (\for_for_j_sva(12)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62989z1419.INIT = 8'h69;
    LUT3 ix62990z1419 (.O (nx62990z2), .I0 (\for_for_j_sva(13)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62990z1419.INIT = 8'h69;
    LUT3 ix62991z1419 (.O (nx62991z2), .I0 (\for_for_j_sva(14)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62991z1419.INIT = 8'h69;
    LUT3 ix62992z1419 (.O (nx62992z2), .I0 (\for_for_j_sva(15)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62992z1419.INIT = 8'h69;
    LUT3 ix62993z1419 (.O (nx62993z2), .I0 (\for_for_j_sva(16)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62993z1419.INIT = 8'h69;
    LUT3 ix62994z1419 (.O (nx62994z2), .I0 (\for_for_j_sva(17)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62994z1419.INIT = 8'h69;
    LUT3 ix62995z1419 (.O (nx62995z2), .I0 (\for_for_j_sva(18)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62995z1419.INIT = 8'h69;
    LUT3 ix62996z1419 (.O (nx62996z2), .I0 (\for_for_j_sva(19)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix62996z1419.INIT = 8'h69;
    LUT3 ix63984z1419 (.O (nx63984z2), .I0 (\for_for_j_sva(20)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63984z1419.INIT = 8'h69;
    LUT3 ix63985z1419 (.O (nx63985z2), .I0 (\for_for_j_sva(21)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63985z1419.INIT = 8'h69;
    LUT3 ix63986z1419 (.O (nx63986z2), .I0 (\for_for_j_sva(22)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63986z1419.INIT = 8'h69;
    LUT3 ix63987z1419 (.O (nx63987z2), .I0 (\for_for_j_sva(23)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63987z1419.INIT = 8'h69;
    LUT3 ix63988z1419 (.O (nx63988z2), .I0 (\for_for_j_sva(24)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63988z1419.INIT = 8'h69;
    LUT3 ix63989z1419 (.O (nx63989z2), .I0 (\for_for_j_sva(25)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63989z1419.INIT = 8'h69;
    LUT3 ix63990z1419 (.O (nx63990z2), .I0 (\for_for_j_sva(26)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63990z1419.INIT = 8'h69;
    LUT3 ix63991z1419 (.O (nx63991z2), .I0 (\for_for_j_sva(27)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63991z1419.INIT = 8'h69;
    LUT3 ix63992z1419 (.O (nx63992z2), .I0 (\for_for_j_sva(28)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63992z1419.INIT = 8'h69;
    LUT3 ix63993z1419 (.O (nx63993z2), .I0 (\for_for_j_sva(29)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63993z1419.INIT = 8'h69;
    LUT3 ix64981z1419 (.O (nx64981z2), .I0 (\for_for_j_sva(30)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix64981z1419.INIT = 8'h69;
    LUT3 ix64982z1419 (.O (nx64982z2), .I0 (\for_for_j_sva(31)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix64982z1419.INIT = 8'h69;
    LUT2 ix8920z1320 (.O (nx8920z1), .I0 (nx12614z3), .I1 (
         conv_core_inst_for_i_sva[31])) ;
         defparam ix8920z1320.INIT = 4'h6;
    LUT2 ix8919z1320 (.O (nx8919z2), .I0 (nx20538z2), .I1 (
         conv_core_inst_for_i_sva[30])) ;
         defparam ix8919z1320.INIT = 4'h6;
    LUT2 ix8918z1320 (.O (nx8918z2), .I0 (nx19541z2), .I1 (
         conv_core_inst_for_i_sva[29])) ;
         defparam ix8918z1320.INIT = 4'h6;
    LUT3 ix8916z1419 (.O (nx8916z2), .I0 (conv_core_inst_for_i_sva[0]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix8916z1419.INIT = 8'h69;
    LUT2 ix34917z1320 (.O (nx34917z1), .I0 (\z_out_4(0)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[12])) ;
         defparam ix34917z1320.INIT = 4'h6;
    LUT2 ix34916z1320 (.O (nx34916z2), .I0 (\z_out_4(1)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[11])) ;
         defparam ix34916z1320.INIT = 4'h6;
    LUT2 ix34915z1320 (.O (nx34915z2), .I0 (\z_out_4(2)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[10])) ;
         defparam ix34915z1320.INIT = 4'h6;
    LUT2 ix34914z1320 (.O (nx34914z2), .I0 (\z_out_4(3)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[9])) ;
         defparam ix34914z1320.INIT = 4'h6;
    LUT2 ix34913z1320 (.O (nx34913z2), .I0 (\z_out_4(4)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[8])) ;
         defparam ix34913z1320.INIT = 4'h6;
    LUT2 ix34912z1320 (.O (nx34912z2), .I0 (\z_out_4(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[7])) ;
         defparam ix34912z1320.INIT = 4'h6;
    LUT2 ix34911z1320 (.O (nx34911z2), .I0 (\z_out_4(6)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[6])) ;
         defparam ix34911z1320.INIT = 4'h6;
    LUT2 ix34910z1320 (.O (nx34910z2), .I0 (\z_out_4(7)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[5])) ;
         defparam ix34910z1320.INIT = 4'h6;
    LUT2 ix34909z1320 (.O (nx34909z2), .I0 (\z_out_4(8)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[4])) ;
         defparam ix34909z1320.INIT = 4'h6;
    LUT2 ix34908z1320 (.O (nx34908z2), .I0 (\z_out_4(9)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[3])) ;
         defparam ix34908z1320.INIT = 4'h6;
    LUT2 ix53948z1320 (.O (nx53948z2), .I0 (\z_out_4(10)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[2])) ;
         defparam ix53948z1320.INIT = 4'h6;
    LUT2 ix53949z1320 (.O (nx53949z2), .I0 (\z_out_4(11)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[1])) ;
         defparam ix53949z1320.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_64" *)
    LUT2 ix38873z1320 (.O (nx38873z2), .I0 (\z_out_4(12)  ), .I1 (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[0])) ;
         defparam ix38873z1320.INIT = 4'h6;
    LUT6 ix28350z14628 (.O (nx28350z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[31]), .I3 (
         conv_core_inst_jj_sva[0]), .I4 (nx28350z4), .I5 (nx28350z5)) ;
         defparam ix28350z14628.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28349z14626 (.O (nx28349z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[30]), .I3 (
         conv_core_inst_jj_sva[1]), .I4 (nx28349z4), .I5 (nx28349z5)) ;
         defparam ix28349z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28348z14626 (.O (nx28348z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[29]), .I3 (
         conv_core_inst_jj_sva[2]), .I4 (nx28348z4), .I5 (nx28348z5)) ;
         defparam ix28348z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28347z14626 (.O (nx28347z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[28]), .I3 (
         conv_core_inst_jj_sva[3]), .I4 (nx28347z4), .I5 (nx28347z5)) ;
         defparam ix28347z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28346z14626 (.O (nx28346z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[27]), .I3 (
         conv_core_inst_jj_sva[4]), .I4 (nx28346z4), .I5 (nx28346z5)) ;
         defparam ix28346z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28345z14626 (.O (nx28345z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[26]), .I3 (
         conv_core_inst_jj_sva[5]), .I4 (nx28345z4), .I5 (nx28345z5)) ;
         defparam ix28345z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28344z14626 (.O (nx28344z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[25]), .I3 (
         conv_core_inst_jj_sva[6]), .I4 (nx28344z4), .I5 (nx28344z5)) ;
         defparam ix28344z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28343z14626 (.O (nx28343z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[24]), .I3 (
         conv_core_inst_jj_sva[7]), .I4 (nx28343z4), .I5 (nx28343z5)) ;
         defparam ix28343z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28342z14626 (.O (nx28342z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[23]), .I3 (
         conv_core_inst_jj_sva[8]), .I4 (nx28342z4), .I5 (nx28342z5)) ;
         defparam ix28342z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix28341z14626 (.O (nx28341z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[22]), .I3 (
         conv_core_inst_jj_sva[9]), .I4 (nx28341z4), .I5 (nx28341z5)) ;
         defparam ix28341z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47647z14626 (.O (nx47647z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[21]), .I3 (
         conv_core_inst_jj_sva[10]), .I4 (nx47647z4), .I5 (nx47647z5)) ;
         defparam ix47647z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47648z14626 (.O (nx47648z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[20]), .I3 (
         conv_core_inst_jj_sva[11]), .I4 (nx47648z4), .I5 (nx47648z5)) ;
         defparam ix47648z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47649z14626 (.O (nx47649z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[19]), .I3 (
         conv_core_inst_jj_sva[12]), .I4 (nx47649z4), .I5 (nx47649z5)) ;
         defparam ix47649z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47650z14626 (.O (nx47650z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[18]), .I3 (
         conv_core_inst_jj_sva[13]), .I4 (nx47650z4), .I5 (nx47650z5)) ;
         defparam ix47650z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47651z14626 (.O (nx47651z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[17]), .I3 (
         conv_core_inst_jj_sva[14]), .I4 (nx47651z4), .I5 (nx47651z5)) ;
         defparam ix47651z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47652z14626 (.O (nx47652z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[16]), .I3 (
         conv_core_inst_jj_sva[15]), .I4 (nx47652z4), .I5 (nx47652z5)) ;
         defparam ix47652z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47653z14626 (.O (nx47653z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[15]), .I3 (
         conv_core_inst_jj_sva[16]), .I4 (nx47653z4), .I5 (nx47653z5)) ;
         defparam ix47653z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47654z14626 (.O (nx47654z4), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[14]), .I3 (
         conv_core_inst_jj_sva[17]), .I4 (nx47654z5), .I5 (nx47654z6)) ;
         defparam ix47654z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47655z14626 (.O (nx47655z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[13]), .I3 (
         conv_core_inst_jj_sva[18]), .I4 (nx47655z4), .I5 (nx47655z5)) ;
         defparam ix47655z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix47656z14626 (.O (nx47656z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[12]), .I3 (
         conv_core_inst_jj_sva[19]), .I4 (nx47656z4), .I5 (nx47656z5)) ;
         defparam ix47656z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48644z14626 (.O (nx48644z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[11]), .I3 (
         conv_core_inst_jj_sva[20]), .I4 (nx48644z4), .I5 (nx48644z5)) ;
         defparam ix48644z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48645z14626 (.O (nx48645z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[10]), .I3 (
         conv_core_inst_jj_sva[21]), .I4 (nx48645z4), .I5 (nx48645z5)) ;
         defparam ix48645z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48646z14626 (.O (nx48646z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[9]), .I3 (
         conv_core_inst_jj_sva[22]), .I4 (nx48646z4), .I5 (nx48646z5)) ;
         defparam ix48646z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48647z14626 (.O (nx48647z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[8]), .I3 (
         conv_core_inst_jj_sva[23]), .I4 (nx48647z4), .I5 (nx48647z5)) ;
         defparam ix48647z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48648z14626 (.O (nx48648z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[7]), .I3 (
         conv_core_inst_jj_sva[24]), .I4 (nx48648z4), .I5 (nx48648z5)) ;
         defparam ix48648z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48649z14626 (.O (nx48649z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[6]), .I3 (
         conv_core_inst_jj_sva[25]), .I4 (nx48649z4), .I5 (nx48649z5)) ;
         defparam ix48649z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48650z14626 (.O (nx48650z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[5]), .I3 (
         conv_core_inst_jj_sva[26]), .I4 (nx48650z4), .I5 (nx48650z5)) ;
         defparam ix48650z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48651z14626 (.O (nx48651z4), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[4]), .I3 (
         conv_core_inst_jj_sva[27]), .I4 (nx48651z5), .I5 (nx48651z6)) ;
         defparam ix48651z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48652z14626 (.O (nx48652z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[3]), .I3 (
         conv_core_inst_jj_sva[28]), .I4 (nx48652z4), .I5 (nx48652z5)) ;
         defparam ix48652z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix48653z14626 (.O (nx48653z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[2]), .I3 (
         conv_core_inst_jj_sva[29]), .I4 (nx48653z4), .I5 (nx48653z5)) ;
         defparam ix48653z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix49641z14626 (.O (nx49641z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(3)  ), .I2 (conv_core_inst_cols_1_sva_1[1]), .I3 (
         conv_core_inst_jj_sva[30]), .I4 (nx49641z4), .I5 (nx49641z5)) ;
         defparam ix49641z14626.INIT = 64'hF1F1C20E000033FF;
    LUT6 ix49642z14524 (.O (nx49642z4), .I0 (nx49642z5), .I1 (\fsm_output(9)  )
         , .I2 (\fsm_output(8)  ), .I3 (nx49642z3), .I4 (
         conv_core_inst_rows_1_sva_2[0]), .I5 (nx49642z6)) ;
         defparam ix49642z14524.INIT = 64'h00AB00ABFF543398;
    INV ix7742z1315 (.O (\kernel_rsci_addr_d_0n0s2(3)  ), .I (
        conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
    INV ix28350z1315 (.O (not_fsm_output_5), .I (\fsm_output(5)  )) ;
    INV ix8917z1315 (.O (\for_for_for_acc_1_psp_sva_11n1s2(3)  ), .I (nx18544z2)
        ) ;
    INV ix62630z1315 (.O (not_fsm_output_4), .I (\fsm_output(4)  )) ;
    (* HLUTNM = "LUT62_1_16" *)
    LUT4 ix49641z14106 (.O (nx49641z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[1]), .I3 (
         \z_out_4(30)  )) ;
         defparam ix49641z14106.INIT = 16'h31F5;
    (* HLUTNM = "LUT62_1_15" *)
    LUT4 ix48653z14106 (.O (nx48653z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[2]), .I3 (
         \z_out_4(29)  )) ;
         defparam ix48653z14106.INIT = 16'h31F5;
    (* HLUTNM = "LUT62_1_14" *)
    LUT4 ix48652z14106 (.O (nx48652z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[3]), .I3 (
         \z_out_4(28)  )) ;
         defparam ix48652z14106.INIT = 16'h31F5;
    (* HLUTNM = "LUT62_1_13" *)
    LUT4 ix48651z14106 (.O (nx48651z6), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[4]), .I3 (
         \z_out_4(27)  )) ;
         defparam ix48651z14106.INIT = 16'h31F5;
    (* HLUTNM = "LUT62_1_12" *)
    LUT4 ix48650z14106 (.O (nx48650z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[5]), .I3 (
         \z_out_4(26)  )) ;
         defparam ix48650z14106.INIT = 16'h31F5;
    (* HLUTNM = "LUT62_1_11" *)
    LUT4 ix48649z14106 (.O (nx48649z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[6]), .I3 (
         \z_out_4(25)  )) ;
         defparam ix48649z14106.INIT = 16'h31F5;
    (* HLUTNM = "LUT62_1_10" *)
    LUT4 ix48648z14106 (.O (nx48648z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[7]), .I3 (
         \z_out_4(24)  )) ;
         defparam ix48648z14106.INIT = 16'h31F5;
    (* HLUTNM = "LUT62_1_9" *)
    LUT4 ix48647z14106 (.O (nx48647z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[8]), .I3 (
         \z_out_4(23)  )) ;
         defparam ix48647z14106.INIT = 16'h31F5;
    LUT4 ix48646z14106 (.O (nx48646z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[9]), .I3 (
         \z_out_4(22)  )) ;
         defparam ix48646z14106.INIT = 16'h31F5;
    LUT4 ix48645z14106 (.O (nx48645z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[10]), .I3 (
         \z_out_4(21)  )) ;
         defparam ix48645z14106.INIT = 16'h31F5;
    LUT4 ix48644z14106 (.O (nx48644z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[11]), .I3 (
         \z_out_4(20)  )) ;
         defparam ix48644z14106.INIT = 16'h31F5;
    LUT4 ix47656z14106 (.O (nx47656z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[12]), .I3 (
         \z_out_4(19)  )) ;
         defparam ix47656z14106.INIT = 16'h31F5;
    LUT4 ix47655z14106 (.O (nx47655z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[13]), .I3 (
         \z_out_4(18)  )) ;
         defparam ix47655z14106.INIT = 16'h31F5;
    LUT4 ix47654z14106 (.O (nx47654z6), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[14]), .I3 (
         conv_core_inst_z_out_4[31])) ;
         defparam ix47654z14106.INIT = 16'h31F5;
    LUT4 ix47653z14106 (.O (nx47653z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[15]), .I3 (
         \z_out_4(16)  )) ;
         defparam ix47653z14106.INIT = 16'h31F5;
    LUT4 ix47652z14106 (.O (nx47652z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[16]), .I3 (
         \z_out_4(15)  )) ;
         defparam ix47652z14106.INIT = 16'h31F5;
    LUT4 ix47651z14106 (.O (nx47651z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[17]), .I3 (
         \z_out_4(14)  )) ;
         defparam ix47651z14106.INIT = 16'h31F5;
    LUT4 ix47650z14106 (.O (nx47650z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[18]), .I3 (
         \z_out_4(13)  )) ;
         defparam ix47650z14106.INIT = 16'h31F5;
    LUT4 ix47649z14106 (.O (nx47649z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[19]), .I3 (
         \z_out_4(12)  )) ;
         defparam ix47649z14106.INIT = 16'h31F5;
    LUT4 ix47648z14106 (.O (nx47648z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[20]), .I3 (
         \z_out_4(11)  )) ;
         defparam ix47648z14106.INIT = 16'h31F5;
    LUT4 ix47647z14106 (.O (nx47647z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[21]), .I3 (
         \z_out_4(10)  )) ;
         defparam ix47647z14106.INIT = 16'h31F5;
    LUT4 ix28341z14106 (.O (nx28341z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[22]), .I3 (
         \z_out_4(9)  )) ;
         defparam ix28341z14106.INIT = 16'h31F5;
    LUT4 ix28342z14106 (.O (nx28342z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[23]), .I3 (
         \z_out_4(8)  )) ;
         defparam ix28342z14106.INIT = 16'h31F5;
    LUT4 ix28343z14106 (.O (nx28343z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[24]), .I3 (
         \z_out_4(7)  )) ;
         defparam ix28343z14106.INIT = 16'h31F5;
    LUT4 ix28344z14106 (.O (nx28344z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[25]), .I3 (
         \z_out_4(6)  )) ;
         defparam ix28344z14106.INIT = 16'h31F5;
    LUT4 ix28345z14106 (.O (nx28345z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[26]), .I3 (
         \z_out_4(5)  )) ;
         defparam ix28345z14106.INIT = 16'h31F5;
    LUT4 ix28346z14106 (.O (nx28346z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[27]), .I3 (
         \z_out_4(4)  )) ;
         defparam ix28346z14106.INIT = 16'h31F5;
    LUT4 ix28347z14106 (.O (nx28347z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[28]), .I3 (
         \z_out_4(3)  )) ;
         defparam ix28347z14106.INIT = 16'h31F5;
    LUT4 ix28348z14106 (.O (nx28348z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[29]), .I3 (
         \z_out_4(2)  )) ;
         defparam ix28348z14106.INIT = 16'h31F5;
    LUT4 ix28349z14106 (.O (nx28349z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[30]), .I3 (
         \z_out_4(1)  )) ;
         defparam ix28349z14106.INIT = 16'h31F5;
    LUT4 ix28350z14108 (.O (nx28350z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_rows_1_sva_2[31]), .I3 (
         \z_out_4(0)  )) ;
         defparam ix28350z14108.INIT = 16'h31F5;
    (* HLUTNM = "LUT62_1_73" *)
    LUT2 ix58321z1320 (.O (nx58321z1), .I0 (nx20538z2), .I1 (nx12614z3)) ;
         defparam ix58321z1320.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_38" *)
    LUT3 ix57324z1400 (.O (nx57324z1), .I0 (nx19541z2), .I1 (nx20538z2), .I2 (
         nx12614z3)) ;
         defparam ix57324z1400.INIT = 8'h56;
    (* HLUTNM = "LUT62_1_1" *)
    LUT4 ix56327z23160 (.O (nx56327z1), .I0 (nx18544z2), .I1 (nx19541z2), .I2 (
         nx20538z2), .I3 (nx12614z3)) ;
         defparam ix56327z23160.INIT = 16'h5556;
    (* HLUTNM = "LUT62_1_1" *)
    LUT5 ix55330z45003 (.O (nx55330z1), .I0 (nx20393z3), .I1 (nx18544z2), .I2 (
         nx19541z2), .I3 (nx20538z2), .I4 (nx12614z3)) ;
         defparam ix55330z45003.INIT = 32'hAAAAAAA9;
    (* HLUTNM = "LUT62_1_17" *)
    LUT4 ix59318z1315 (.O (nx59318z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  )) ;
         defparam ix59318z1315.INIT = 16'h0001;
    (* HLUTNM = "LUT62_1_7" *)
    LUT4 ix21003z3405 (.O (nx21003z2), .I0 (\fsm_output(7)  ), .I1 (
         \fsm_output(3)  ), .I2 (\for_for_for_for_n_4_0_sva(0)  ), .I3 (
         nx12614z3)) ;
         defparam ix21003z3405.INIT = 16'h082A;
    LUT6 ix22000z3490 (.O (nx22000z1), .I0 (\fsm_output(7)  ), .I1 (
         \fsm_output(3)  ), .I2 (\for_for_for_for_n_4_0_sva(1)  ), .I3 (
         \for_for_for_for_n_4_0_sva(0)  ), .I4 (nx20538z2), .I5 (nx12614z3)) ;
         defparam ix22000z3490.INIT = 64'h08802AA22AA20880;
    LUT6 ix22997z42914 (.O (nx22997z1), .I0 (\fsm_output(7)  ), .I1 (
         \fsm_output(3)  ), .I2 (\for_for_for_for_n_4_0_sva(2)  ), .I3 (
         nx19541z2), .I4 (nx12614z2), .I5 (nx20393z4)) ;
         defparam ix22997z42914.INIT = 64'hA280082AA280A280;
    (* HLUTNM = "LUT62_1_7" *)
    LUT2 ix23994z1322 (.O (nx23994z1), .I0 (\fsm_output(7)  ), .I1 (nx18544z1)
         ) ;
         defparam ix23994z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_63" *)
    LUT2 ix24991z1322 (.O (nx24991z1), .I0 (\fsm_output(7)  ), .I1 (nx20393z2)
         ) ;
         defparam ix24991z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_4" *)
    LUT3 ix21003z1568 (.O (nx21003z1), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(7)  ), .I2 (\fsm_output(1)  )) ;
         defparam ix21003z1568.INIT = 8'hFE;
    (* HLUTNM = "LUT62_1_5" *)
    LUT3 ix15408z1562 (.O (nx15408z1), .I0 (\fsm_output(6)  ), .I1 (
         for_for_for_for_slc_for_for_for_for_acc_5_itm), .I2 (
         \conv_core_core_fsm_inst_fsm_output(2)  )) ;
         defparam ix15408z1562.INIT = 8'hF8;
    (* HLUTNM = "LUT62_1_5" *)
    LUT2 ix19396z1316 (.O (nx19396z1), .I0 (\fsm_output(6)  ), .I1 (
         for_for_for_for_slc_for_for_for_for_acc_5_itm)) ;
         defparam ix19396z1316.INIT = 4'h2;
    LUT6 ix20393z42404 (.O (nx20393z1), .I0 (\fsm_output(7)  ), .I1 (nx12614z2)
         , .I2 (nx20393z2), .I3 (nx18544z1), .I4 (nx19541z1), .I5 (nx20538z1)) ;
         defparam ix20393z42404.INIT = 64'hA0A0A0A0A0A0A082;
    (* HLUTNM = "LUT62_1_65" *)
    LUT2 ix43133z1328 (.O (nx43133z1), .I0 (p_rst_int), .I1 (\p_fsm_output(10)  
         )) ;
         defparam ix43133z1328.INIT = 4'hE;
    LUT5 ix60570z1316 (.O (nx60570z1), .I0 (\z_out_1(32)  ), .I1 (nx60570z2), .I2 (
         conv_core_inst_jj_sva[31]), .I3 (
         conv_core_inst_for_for_for_for_acc_3_tmp[31]), .I4 (
         conv_core_inst_rows_1_sva_2[0])) ;
         defparam ix60570z1316.INIT = 32'h00000002;
    LUT5 ix12614z14424 (.O (nx12614z1), .I0 (nx12614z2), .I1 (nx20393z2), .I2 (
         nx18544z1), .I3 (nx19541z1), .I4 (nx20538z1)) ;
         defparam ix12614z14424.INIT = 32'h33333336;
    (* HLUTNM = "LUT62_1_3" *)
    LUT5 ix20538z33354 (.O (nx20538z1), .I0 (\fsm_output(3)  ), .I1 (
         \for_for_for_for_n_4_0_sva(1)  ), .I2 (\for_for_for_for_n_4_0_sva(0)  )
         , .I3 (nx20538z2), .I4 (nx12614z3)) ;
         defparam ix20538z33354.INIT = 32'h287D7D28;
    LUT6 ix19541z33354 (.O (nx19541z1), .I0 (\fsm_output(3)  ), .I1 (
         \for_for_for_for_n_4_0_sva(2)  ), .I2 (\for_for_for_for_n_4_0_sva(1)  )
         , .I3 (nx19541z2), .I4 (nx20538z2), .I5 (nx12614z2)) ;
         defparam ix19541z33354.INIT = 64'hDD88DD88287D7D28;
    LUT6 ix18544z56826 (.O (nx18544z1), .I0 (\fsm_output(3)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4]), .I2 (nx18544z2), .I3 (
         nx12614z2), .I4 (nx20393z4), .I5 (nx18544z3)) ;
         defparam ix18544z56826.INIT = 64'hD827D8D8D8D8D8D8;
    (* HLUTNM = "LUT62_1_2" *)
    LUT3 ix18544z1531 (.O (nx18544z3), .I0 (\fsm_output(3)  ), .I1 (
         \for_for_for_for_n_4_0_sva(2)  ), .I2 (nx19541z2)) ;
         defparam ix18544z1531.INIT = 8'hD8;
    LUT6 ix20393z56827 (.O (nx20393z2), .I0 (\fsm_output(3)  ), .I1 (
         \for_for_for_for_n_4_0_sva(4)  ), .I2 (nx20393z3), .I3 (nx12614z2), .I4 (
         nx20393z4), .I5 (nx20393z5)) ;
         defparam ix20393z56827.INIT = 64'hD827D8D8D8D8D8D8;
    (* HLUTNM = "LUT62_1_2" *)
    LUT5 ix20393z34213 (.O (nx20393z5), .I0 (\fsm_output(3)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4]), .I2 (
         \for_for_for_for_n_4_0_sva(2)  ), .I3 (nx18544z2), .I4 (nx19541z2)) ;
         defparam ix20393z34213.INIT = 32'hD5808080;
    (* HLUTNM = "LUT62_1_38" *)
    LUT3 ix20393z1532 (.O (nx20393z4), .I0 (\fsm_output(3)  ), .I1 (
         \for_for_for_for_n_4_0_sva(1)  ), .I2 (nx20538z2)) ;
         defparam ix20393z1532.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_3" *)
    LUT3 ix12614z1354 (.O (nx12614z2), .I0 (\fsm_output(3)  ), .I1 (
         \for_for_for_for_n_4_0_sva(0)  ), .I2 (nx12614z3)) ;
         defparam ix12614z1354.INIT = 8'h27;
    (* HLUTNM = "LUT62_1_29" *)
    LUT2 ix33183z1322 (.O (nx33183z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(0)  
         )) ;
         defparam ix33183z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_27" *)
    LUT2 ix32186z1322 (.O (nx32186z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(1)  
         )) ;
         defparam ix32186z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_25" *)
    LUT2 ix31189z1322 (.O (nx31189z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(2)  
         )) ;
         defparam ix31189z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_23" *)
    LUT2 ix30192z1322 (.O (nx30192z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(3)  
         )) ;
         defparam ix30192z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_22" *)
    LUT2 ix29195z1322 (.O (nx29195z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(4)  
         )) ;
         defparam ix29195z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_21" *)
    LUT2 ix28198z1322 (.O (nx28198z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(5)  
         )) ;
         defparam ix28198z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_20" *)
    LUT2 ix27201z1322 (.O (nx27201z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(6)  
         )) ;
         defparam ix27201z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_19" *)
    LUT2 ix26204z1322 (.O (nx26204z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(7)  
         )) ;
         defparam ix26204z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_18" *)
    LUT2 ix25207z1322 (.O (nx25207z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(8)  
         )) ;
         defparam ix25207z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_6" *)
    LUT2 ix24210z1322 (.O (nx24210z1), .I0 (\fsm_output(8)  ), .I1 (\z_out_2(9)  
         )) ;
         defparam ix24210z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_24" *)
    LUT2 ix30218z1322 (.O (nx30218z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(10)  )) ;
         defparam ix30218z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_26" *)
    LUT2 ix31215z1322 (.O (nx31215z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(11)  )) ;
         defparam ix31215z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_28" *)
    LUT2 ix32212z1322 (.O (nx32212z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(12)  )) ;
         defparam ix32212z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_30" *)
    LUT2 ix33209z1322 (.O (nx33209z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(13)  )) ;
         defparam ix33209z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_31" *)
    LUT2 ix34206z1322 (.O (nx34206z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(14)  )) ;
         defparam ix34206z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_32" *)
    LUT2 ix35203z1322 (.O (nx35203z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(15)  )) ;
         defparam ix35203z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_33" *)
    LUT2 ix36200z1322 (.O (nx36200z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(16)  )) ;
         defparam ix36200z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_34" *)
    LUT2 ix37197z1322 (.O (nx37197z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(17)  )) ;
         defparam ix37197z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_35" *)
    LUT2 ix38194z1322 (.O (nx38194z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(18)  )) ;
         defparam ix38194z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_36" *)
    LUT2 ix39191z1322 (.O (nx39191z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(19)  )) ;
         defparam ix39191z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_37" *)
    LUT2 ix41187z1322 (.O (nx41187z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(20)  )) ;
         defparam ix41187z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_64" *)
    LUT2 ix42184z1322 (.O (nx42184z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(21)  )) ;
         defparam ix42184z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_65" *)
    LUT2 ix43181z1322 (.O (nx43181z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(22)  )) ;
         defparam ix43181z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_47" *)
    LUT2 ix44178z1322 (.O (nx44178z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(23)  )) ;
         defparam ix44178z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_47" *)
    LUT2 ix45175z1322 (.O (nx45175z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(24)  )) ;
         defparam ix45175z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_66" *)
    LUT2 ix46172z1322 (.O (nx46172z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(25)  )) ;
         defparam ix46172z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_68" *)
    LUT2 ix47169z1322 (.O (nx47169z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(26)  )) ;
         defparam ix47169z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_69" *)
    LUT2 ix48166z1322 (.O (nx48166z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(27)  )) ;
         defparam ix48166z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_70" *)
    LUT2 ix49163z1322 (.O (nx49163z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(28)  )) ;
         defparam ix49163z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_71" *)
    LUT2 ix50160z1322 (.O (nx50160z1), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(29)  )) ;
         defparam ix50160z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_51" *)
    LUT2 ix52156z1323 (.O (nx52156z2), .I0 (\fsm_output(8)  ), .I1 (
         \z_out_2(30)  )) ;
         defparam ix52156z1323.INIT = 4'h8;
    LUT6 ix53153z53742 (.O (nx53153z1), .I0 (p_nbus_rows_rsc_z_int[0]), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(0)  ), .I3 (\for_for_j_sva(31)  ), 
         .I4 (nx21390z2), .I5 (nx22387z2)) ;
         defparam ix53153z53742.INIT = 64'h008CCC400000CCCC;
    (* HLUTNM = "LUT62_1_51" *)
    LUT2 ix52156z1328 (.O (nx52156z1), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  )) ;
         defparam ix52156z1328.INIT = 4'hE;
    (* HLUTNM = "LUT62_1_50" *)
    LUT2 ix51642z1322 (.O (nx51642z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(0)  
         )) ;
         defparam ix51642z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_49" *)
    LUT2 ix50645z1322 (.O (nx50645z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(1)  
         )) ;
         defparam ix50645z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_71" *)
    LUT2 ix49648z1322 (.O (nx49648z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(2)  
         )) ;
         defparam ix49648z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_48" *)
    LUT2 ix48651z1322 (.O (nx48651z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(3)  
         )) ;
         defparam ix48651z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_69" *)
    LUT2 ix47654z1322 (.O (nx47654z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(4)  
         )) ;
         defparam ix47654z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_67" *)
    LUT2 ix46657z1322 (.O (nx46657z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(5)  
         )) ;
         defparam ix46657z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_16" *)
    LUT2 ix45660z1322 (.O (nx45660z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(6)  
         )) ;
         defparam ix45660z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_14" *)
    LUT2 ix44663z1322 (.O (nx44663z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(7)  
         )) ;
         defparam ix44663z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_12" *)
    LUT2 ix43666z1322 (.O (nx43666z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(8)  
         )) ;
         defparam ix43666z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_10" *)
    LUT2 ix42669z1322 (.O (nx42669z1), .I0 (\fsm_output(9)  ), .I1 (\z_out_2(9)  
         )) ;
         defparam ix42669z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_8" *)
    LUT2 ix42211z1322 (.O (nx42211z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(10)  )) ;
         defparam ix42211z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_11" *)
    LUT2 ix43208z1322 (.O (nx43208z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(11)  )) ;
         defparam ix43208z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_13" *)
    LUT2 ix44205z1322 (.O (nx44205z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(12)  )) ;
         defparam ix44205z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_15" *)
    LUT2 ix45202z1322 (.O (nx45202z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(13)  )) ;
         defparam ix45202z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_66" *)
    LUT2 ix46199z1322 (.O (nx46199z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(14)  )) ;
         defparam ix46199z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_68" *)
    LUT2 ix47196z1322 (.O (nx47196z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(15)  )) ;
         defparam ix47196z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_48" *)
    LUT2 ix48193z1322 (.O (nx48193z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(16)  )) ;
         defparam ix48193z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_70" *)
    LUT2 ix49190z1322 (.O (nx49190z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(17)  )) ;
         defparam ix49190z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_49" *)
    LUT2 ix50187z1322 (.O (nx50187z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(18)  )) ;
         defparam ix50187z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_50" *)
    LUT2 ix51184z1322 (.O (nx51184z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(19)  )) ;
         defparam ix51184z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_52" *)
    LUT2 ix53180z1322 (.O (nx53180z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(20)  )) ;
         defparam ix53180z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_52" *)
    LUT2 ix54177z1322 (.O (nx54177z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(21)  )) ;
         defparam ix54177z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_53" *)
    LUT2 ix55174z1322 (.O (nx55174z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(22)  )) ;
         defparam ix55174z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_53" *)
    LUT2 ix56171z1322 (.O (nx56171z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(23)  )) ;
         defparam ix56171z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_72" *)
    LUT2 ix57168z1322 (.O (nx57168z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(24)  )) ;
         defparam ix57168z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_73" *)
    LUT2 ix58165z1322 (.O (nx58165z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(25)  )) ;
         defparam ix58165z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_54" *)
    LUT2 ix59162z1322 (.O (nx59162z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(26)  )) ;
         defparam ix59162z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_54" *)
    LUT2 ix60159z1322 (.O (nx60159z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(27)  )) ;
         defparam ix60159z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_55" *)
    LUT2 ix61156z1322 (.O (nx61156z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(28)  )) ;
         defparam ix61156z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_55" *)
    LUT2 ix62153z1322 (.O (nx62153z1), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(29)  )) ;
         defparam ix62153z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_74" *)
    LUT2 ix64149z1323 (.O (nx64149z2), .I0 (\fsm_output(9)  ), .I1 (
         \z_out_2(30)  )) ;
         defparam ix64149z1323.INIT = 4'h8;
    LUT6 ix65146z45004 (.O (nx65146z1), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[0]), .I3 (
         conv_core_inst_for_i_sva[27]), .I4 (nx21390z2), .I5 (nx13414z2)) ;
         defparam ix65146z45004.INIT = 64'h00A2AA080000AAAA;
    LUT2 ix64149z1328 (.O (nx64149z1), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(0)  )) ;
         defparam ix64149z1328.INIT = 4'hE;
    LUT2 ix9631z1328 (.O (nx9631z1), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(0)  )) ;
         defparam ix9631z1328.INIT = 4'hE;
    (* HLUTNM = "LUT62_1_72" *)
    LUT2 ix5701z1322 (.O (nx5701z1), .I0 (\fsm_output(6)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[4])) ;
         defparam ix5701z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_67" *)
    LUT2 ix4704z1322 (.O (nx4704z1), .I0 (\fsm_output(6)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[3])) ;
         defparam ix4704z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_46" *)
    LUT2 ix3707z1322 (.O (nx3707z1), .I0 (\fsm_output(6)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[2])) ;
         defparam ix3707z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_46" *)
    LUT2 ix2710z1322 (.O (nx2710z1), .I0 (\fsm_output(6)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[1])) ;
         defparam ix2710z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_17" *)
    LUT2 ix1713z1322 (.O (nx1713z1), .I0 (\fsm_output(6)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva_3[0])) ;
         defparam ix1713z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_74" *)
    LUT2 ix63825z1336 (.O (nx63825z15), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[14])) ;
         defparam ix63825z1336.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_62" *)
    LUT2 ix63825z1335 (.O (nx63825z14), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[13])) ;
         defparam ix63825z1335.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_62" *)
    LUT2 ix63825z1334 (.O (nx63825z13), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[12])) ;
         defparam ix63825z1334.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_61" *)
    LUT2 ix63825z1333 (.O (nx63825z12), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[11])) ;
         defparam ix63825z1333.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_61" *)
    LUT2 ix63825z1332 (.O (nx63825z11), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[10])) ;
         defparam ix63825z1332.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_60" *)
    LUT2 ix63825z1331 (.O (nx63825z10), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[9])) ;
         defparam ix63825z1331.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_60" *)
    LUT2 ix63825z1330 (.O (nx63825z9), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[8])) ;
         defparam ix63825z1330.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_59" *)
    LUT2 ix63825z1329 (.O (nx63825z8), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[7])) ;
         defparam ix63825z1329.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_59" *)
    LUT2 ix63825z1328 (.O (nx63825z7), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[6])) ;
         defparam ix63825z1328.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_58" *)
    LUT2 ix63825z1327 (.O (nx63825z6), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[5])) ;
         defparam ix63825z1327.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_58" *)
    LUT2 ix63825z1326 (.O (nx63825z5), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[4])) ;
         defparam ix63825z1326.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_57" *)
    LUT2 ix63825z1325 (.O (nx63825z4), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[3])) ;
         defparam ix63825z1325.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_57" *)
    LUT2 ix63825z1324 (.O (nx63825z3), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[2])) ;
         defparam ix63825z1324.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_56" *)
    LUT2 ix63825z1323 (.O (nx63825z2), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[1])) ;
         defparam ix63825z1323.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_56" *)
    LUT2 ix63825z1322 (.O (nx63825z1), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[0])) ;
         defparam ix63825z1322.INIT = 4'h8;
    LUT4 ix18281z64952 (.O (nx18281z15), .I0 (p_nbus_image_rsc_data_out_int[0])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64952.INIT = 16'hF888;
    LUT4 ix18281z64951 (.O (nx18281z14), .I0 (p_nbus_image_rsc_data_out_int[1])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64951.INIT = 16'hF888;
    LUT4 ix18281z64950 (.O (nx18281z13), .I0 (p_nbus_image_rsc_data_out_int[2])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64950.INIT = 16'hF888;
    LUT4 ix18281z64949 (.O (nx18281z12), .I0 (p_nbus_image_rsc_data_out_int[3])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64949.INIT = 16'hF888;
    LUT4 ix18281z64948 (.O (nx18281z11), .I0 (p_nbus_image_rsc_data_out_int[4])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64948.INIT = 16'hF888;
    LUT4 ix18281z64947 (.O (nx18281z10), .I0 (p_nbus_image_rsc_data_out_int[5])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64947.INIT = 16'hF888;
    LUT4 ix18281z64946 (.O (nx18281z9), .I0 (p_nbus_image_rsc_data_out_int[6]), 
         .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64946.INIT = 16'hF888;
    LUT4 ix18281z64945 (.O (nx18281z8), .I0 (p_nbus_image_rsc_data_out_int[7]), 
         .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64945.INIT = 16'hF888;
    LUT4 ix18281z64944 (.O (nx18281z7), .I0 (p_nbus_image_rsc_data_out_int[8]), 
         .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64944.INIT = 16'hF888;
    LUT4 ix18281z64943 (.O (nx18281z6), .I0 (p_nbus_image_rsc_data_out_int[9]), 
         .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64943.INIT = 16'hF888;
    LUT4 ix18281z64942 (.O (nx18281z5), .I0 (p_nbus_image_rsc_data_out_int[10])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64942.INIT = 16'hF888;
    LUT4 ix18281z64941 (.O (nx18281z4), .I0 (p_nbus_image_rsc_data_out_int[11])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64941.INIT = 16'hF888;
    LUT4 ix18281z64940 (.O (nx18281z3), .I0 (p_nbus_image_rsc_data_out_int[12])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64940.INIT = 16'hF888;
    LUT4 ix18281z64939 (.O (nx18281z2), .I0 (p_nbus_image_rsc_data_out_int[13])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64939.INIT = 16'hF888;
    LUT4 ix18281z64938 (.O (nx18281z1), .I0 (p_nbus_image_rsc_data_out_int[14])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix18281z64938.INIT = 16'hF888;
    LUT4 ix30685z1087 (.O (nx30685z34), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(4)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[31])) ;
         defparam ix30685z1087.INIT = 16'hFEFC;
    LUT3 ix30685z1582 (.O (nx30685z33), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[30])) ;
         defparam ix30685z1582.INIT = 8'hEC;
    LUT2 ix30685z1353 (.O (nx30685z32), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[29])) ;
         defparam ix30685z1353.INIT = 4'h8;
    LUT4 ix30685z1084 (.O (nx30685z31), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(4)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[28])) ;
         defparam ix30685z1084.INIT = 16'hFEFC;
    LUT4 ix30685z1083 (.O (nx30685z30), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(4)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[27])) ;
         defparam ix30685z1083.INIT = 16'hFEFC;
    LUT2 ix30685z1350 (.O (nx30685z29), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[26])) ;
         defparam ix30685z1350.INIT = 4'h8;
    LUT2 ix30685z1349 (.O (nx30685z28), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[25])) ;
         defparam ix30685z1349.INIT = 4'h8;
    LUT2 ix30685z1348 (.O (nx30685z27), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[24])) ;
         defparam ix30685z1348.INIT = 4'h8;
    LUT2 ix30685z1347 (.O (nx30685z26), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[23])) ;
         defparam ix30685z1347.INIT = 4'h8;
    LUT2 ix30685z1346 (.O (nx30685z25), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[22])) ;
         defparam ix30685z1346.INIT = 4'h8;
    LUT2 ix30685z1345 (.O (nx30685z24), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[21])) ;
         defparam ix30685z1345.INIT = 4'h8;
    LUT2 ix30685z1344 (.O (nx30685z23), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[20])) ;
         defparam ix30685z1344.INIT = 4'h8;
    LUT2 ix30685z1343 (.O (nx30685z22), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[19])) ;
         defparam ix30685z1343.INIT = 4'h8;
    LUT2 ix30685z1342 (.O (nx30685z21), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[18])) ;
         defparam ix30685z1342.INIT = 4'h8;
    LUT2 ix30685z1341 (.O (nx30685z20), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[17])) ;
         defparam ix30685z1341.INIT = 4'h8;
    LUT2 ix30685z1340 (.O (nx30685z19), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[16])) ;
         defparam ix30685z1340.INIT = 4'h8;
    LUT2 ix30685z1339 (.O (nx30685z18), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[15])) ;
         defparam ix30685z1339.INIT = 4'h8;
    LUT6 ix30685z36282 (.O (nx30685z17), .I0 (p_nbus_image_rsc_data_out_int[15])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[31]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[12])) ;
         defparam ix30685z36282.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36281 (.O (nx30685z16), .I0 (p_nbus_image_rsc_data_out_int[16])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[30]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[11])) ;
         defparam ix30685z36281.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36280 (.O (nx30685z15), .I0 (p_nbus_image_rsc_data_out_int[17])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[29]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[10])) ;
         defparam ix30685z36280.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36279 (.O (nx30685z14), .I0 (p_nbus_image_rsc_data_out_int[18])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[28]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[9])) ;
         defparam ix30685z36279.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36278 (.O (nx30685z13), .I0 (p_nbus_image_rsc_data_out_int[19])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[0]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[8])) ;
         defparam ix30685z36278.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36277 (.O (nx30685z12), .I0 (p_nbus_image_rsc_data_out_int[20])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[1]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[7])) ;
         defparam ix30685z36277.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36276 (.O (nx30685z11), .I0 (p_nbus_image_rsc_data_out_int[21])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[2]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[6])) ;
         defparam ix30685z36276.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36275 (.O (nx30685z10), .I0 (p_nbus_image_rsc_data_out_int[22])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[3]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[5])) ;
         defparam ix30685z36275.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36274 (.O (nx30685z9), .I0 (p_nbus_image_rsc_data_out_int[23])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[4]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[4])) ;
         defparam ix30685z36274.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36273 (.O (nx30685z8), .I0 (p_nbus_image_rsc_data_out_int[24])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[5]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[3])) ;
         defparam ix30685z36273.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36272 (.O (nx30685z7), .I0 (p_nbus_image_rsc_data_out_int[25])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[6]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[2])) ;
         defparam ix30685z36272.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36271 (.O (nx30685z6), .I0 (p_nbus_image_rsc_data_out_int[26])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[7]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[1])) ;
         defparam ix30685z36271.INIT = 64'hFFF8F8F8FF888888;
    LUT6 ix30685z36270 (.O (nx30685z5), .I0 (p_nbus_image_rsc_data_out_int[27])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(4)  ), .I3 (\fsm_output(3)  
         ), .I4 (conv_core_inst_for_i_sva[8]), .I5 (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[0])) ;
         defparam ix30685z36270.INIT = 64'hFFF8F8F8FF888888;
    LUT4 ix30685z64941 (.O (nx30685z4), .I0 (p_nbus_image_rsc_data_out_int[28])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix30685z64941.INIT = 16'hF888;
    LUT4 ix30685z64940 (.O (nx30685z3), .I0 (p_nbus_image_rsc_data_out_int[29])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix30685z64940.INIT = 16'hF888;
    LUT4 ix30685z64939 (.O (nx30685z2), .I0 (p_nbus_image_rsc_data_out_int[30])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix30685z64939.INIT = 16'hF888;
    LUT4 ix30685z64938 (.O (nx30685z1), .I0 (p_nbus_image_rsc_data_out_int[31])
         , .I1 (\fsm_output(5)  ), .I2 (\fsm_output(3)  ), .I3 (
         conv_core_inst_for_i_sva[9])) ;
         defparam ix30685z64938.INIT = 16'hF888;
    LUT6 ix49642z4912 (.O (nx49642z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (nx21390z2), .I3 (nx22387z2), .I4 (nx13414z2), .I5 (
         nx49642z3)) ;
         defparam ix49642z4912.INIT = 64'hFFFFFFFFE00E0E0E;
    LUT6 ix49642z1317 (.O (nx49642z5), .I0 (\fsm_output(9)  ), .I1 (
         conv_core_inst_cols_1_sva_1[0]), .I2 (\fsm_output(1)  ), .I3 (
         conv_core_inst_for_i_sva[27]), .I4 (nx21390z2), .I5 (nx13414z2)) ;
         defparam ix49642z1317.INIT = 64'hBA3045CFFFFF0000;
    LUT6 ix14411z1314 (.O (nx14411z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[0]), .I3 (
         conv_core_inst_for_i_sva[27]), .I4 (nx21390z2), .I5 (nx13414z2)) ;
         defparam ix14411z1314.INIT = 64'h0000AE0C0000FFFF;
    LUT4 ix49642z61891 (.O (nx49642z3), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[0]), .I3 (
         conv_core_inst_jj_sva[31])) ;
         defparam ix49642z61891.INIT = 16'hECA0;
    (* HLUTNM = "LUT62_1_6" *)
    LUT4 ix13414z10450 (.O (nx13414z2), .I0 (p_nbus_rows_rsc_z_int[0]), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(0)  ), .I3 (\for_for_j_sva(31)  )
         ) ;
         defparam ix13414z10450.INIT = 16'h23AF;
    (* HLUTNM = "LUT62_1_8" *)
    LUT4 ix22387z22294 (.O (nx22387z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[0]), .I3 (
         conv_core_inst_for_i_sva[27])) ;
         defparam ix22387z22294.INIT = 16'h51F3;
    LUT6 ix49641z61890 (.O (nx49641z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[1]), .I3 (
         conv_core_inst_jj_sva[30]), .I4 (\z_out_2(30)  ), .I5 (nx28350z2)) ;
         defparam ix49641z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix49641z62756 (.O (nx49641z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[1]), .I4 (\z_out_2(30)  )
         ) ;
         defparam ix49641z62756.INIT = 32'hFEEEF000;
    LUT6 ix48653z61890 (.O (nx48653z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[2]), .I3 (
         conv_core_inst_jj_sva[29]), .I4 (\z_out_2(29)  ), .I5 (nx28350z2)) ;
         defparam ix48653z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48653z62756 (.O (nx48653z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[2]), .I4 (\z_out_2(29)  )
         ) ;
         defparam ix48653z62756.INIT = 32'hFEEEF000;
    LUT6 ix48652z61890 (.O (nx48652z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[3]), .I3 (
         conv_core_inst_jj_sva[28]), .I4 (\z_out_2(28)  ), .I5 (nx28350z2)) ;
         defparam ix48652z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48652z62756 (.O (nx48652z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[3]), .I4 (\z_out_2(28)  )
         ) ;
         defparam ix48652z62756.INIT = 32'hFEEEF000;
    LUT6 ix48651z61890 (.O (nx48651z3), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[4]), .I3 (
         conv_core_inst_jj_sva[27]), .I4 (\z_out_2(27)  ), .I5 (nx28350z2)) ;
         defparam ix48651z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48651z62756 (.O (nx48651z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[4]), .I4 (\z_out_2(27)  )
         ) ;
         defparam ix48651z62756.INIT = 32'hFEEEF000;
    LUT6 ix48650z61890 (.O (nx48650z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[5]), .I3 (
         conv_core_inst_jj_sva[26]), .I4 (\z_out_2(26)  ), .I5 (nx28350z2)) ;
         defparam ix48650z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48650z62756 (.O (nx48650z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[5]), .I4 (\z_out_2(26)  )
         ) ;
         defparam ix48650z62756.INIT = 32'hFEEEF000;
    LUT6 ix48649z61890 (.O (nx48649z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[6]), .I3 (
         conv_core_inst_jj_sva[25]), .I4 (\z_out_2(25)  ), .I5 (nx28350z2)) ;
         defparam ix48649z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48649z62756 (.O (nx48649z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[6]), .I4 (\z_out_2(25)  )
         ) ;
         defparam ix48649z62756.INIT = 32'hFEEEF000;
    LUT6 ix48648z61890 (.O (nx48648z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[7]), .I3 (
         conv_core_inst_jj_sva[24]), .I4 (\z_out_2(24)  ), .I5 (nx28350z2)) ;
         defparam ix48648z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48648z62756 (.O (nx48648z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[7]), .I4 (\z_out_2(24)  )
         ) ;
         defparam ix48648z62756.INIT = 32'hFEEEF000;
    LUT6 ix48647z61890 (.O (nx48647z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[8]), .I3 (
         conv_core_inst_jj_sva[23]), .I4 (\z_out_2(23)  ), .I5 (nx28350z2)) ;
         defparam ix48647z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48647z62756 (.O (nx48647z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[8]), .I4 (\z_out_2(23)  )
         ) ;
         defparam ix48647z62756.INIT = 32'hFEEEF000;
    LUT6 ix48646z61890 (.O (nx48646z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[9]), .I3 (
         conv_core_inst_jj_sva[22]), .I4 (\z_out_2(22)  ), .I5 (nx28350z2)) ;
         defparam ix48646z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48646z62756 (.O (nx48646z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[9]), .I4 (\z_out_2(22)  )
         ) ;
         defparam ix48646z62756.INIT = 32'hFEEEF000;
    LUT6 ix48645z61890 (.O (nx48645z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[10]), .I3 (
         conv_core_inst_jj_sva[21]), .I4 (\z_out_2(21)  ), .I5 (nx28350z2)) ;
         defparam ix48645z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48645z62756 (.O (nx48645z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[10]), .I4 (\z_out_2(21)  
         )) ;
         defparam ix48645z62756.INIT = 32'hFEEEF000;
    LUT6 ix48644z61890 (.O (nx48644z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[11]), .I3 (
         conv_core_inst_jj_sva[20]), .I4 (\z_out_2(20)  ), .I5 (nx28350z2)) ;
         defparam ix48644z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix48644z62756 (.O (nx48644z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[11]), .I4 (\z_out_2(20)  
         )) ;
         defparam ix48644z62756.INIT = 32'hFEEEF000;
    LUT6 ix47656z61890 (.O (nx47656z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[12]), .I3 (
         conv_core_inst_jj_sva[19]), .I4 (\z_out_2(19)  ), .I5 (nx28350z2)) ;
         defparam ix47656z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47656z62756 (.O (nx47656z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[12]), .I4 (\z_out_2(19)  
         )) ;
         defparam ix47656z62756.INIT = 32'hFEEEF000;
    LUT6 ix47655z61890 (.O (nx47655z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[13]), .I3 (
         conv_core_inst_jj_sva[18]), .I4 (\z_out_2(18)  ), .I5 (nx28350z2)) ;
         defparam ix47655z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47655z62756 (.O (nx47655z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[13]), .I4 (\z_out_2(18)  
         )) ;
         defparam ix47655z62756.INIT = 32'hFEEEF000;
    LUT6 ix47654z61890 (.O (nx47654z3), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[14]), .I3 (
         conv_core_inst_jj_sva[17]), .I4 (\z_out_2(17)  ), .I5 (nx28350z2)) ;
         defparam ix47654z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47654z62756 (.O (nx47654z5), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[14]), .I4 (\z_out_2(17)  
         )) ;
         defparam ix47654z62756.INIT = 32'hFEEEF000;
    LUT6 ix47653z61890 (.O (nx47653z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[15]), .I3 (
         conv_core_inst_jj_sva[16]), .I4 (\z_out_2(16)  ), .I5 (nx28350z2)) ;
         defparam ix47653z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47653z62756 (.O (nx47653z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[15]), .I4 (\z_out_2(16)  
         )) ;
         defparam ix47653z62756.INIT = 32'hFEEEF000;
    LUT6 ix47652z61890 (.O (nx47652z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[16]), .I3 (
         conv_core_inst_jj_sva[15]), .I4 (\z_out_2(15)  ), .I5 (nx28350z2)) ;
         defparam ix47652z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47652z62756 (.O (nx47652z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[16]), .I4 (\z_out_2(15)  
         )) ;
         defparam ix47652z62756.INIT = 32'hFEEEF000;
    LUT6 ix47651z61890 (.O (nx47651z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[17]), .I3 (
         conv_core_inst_jj_sva[14]), .I4 (\z_out_2(14)  ), .I5 (nx28350z2)) ;
         defparam ix47651z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47651z62756 (.O (nx47651z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[17]), .I4 (\z_out_2(14)  
         )) ;
         defparam ix47651z62756.INIT = 32'hFEEEF000;
    LUT6 ix47650z61890 (.O (nx47650z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[18]), .I3 (
         conv_core_inst_jj_sva[13]), .I4 (\z_out_2(13)  ), .I5 (nx28350z2)) ;
         defparam ix47650z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47650z62756 (.O (nx47650z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[18]), .I4 (\z_out_2(13)  
         )) ;
         defparam ix47650z62756.INIT = 32'hFEEEF000;
    LUT6 ix47649z61890 (.O (nx47649z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[19]), .I3 (
         conv_core_inst_jj_sva[12]), .I4 (\z_out_2(12)  ), .I5 (nx28350z2)) ;
         defparam ix47649z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47649z62756 (.O (nx47649z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[19]), .I4 (\z_out_2(12)  
         )) ;
         defparam ix47649z62756.INIT = 32'hFEEEF000;
    LUT6 ix47648z61890 (.O (nx47648z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[20]), .I3 (
         conv_core_inst_jj_sva[11]), .I4 (\z_out_2(11)  ), .I5 (nx28350z2)) ;
         defparam ix47648z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47648z62756 (.O (nx47648z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[20]), .I4 (\z_out_2(11)  
         )) ;
         defparam ix47648z62756.INIT = 32'hFEEEF000;
    LUT6 ix47647z61890 (.O (nx47647z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[21]), .I3 (
         conv_core_inst_jj_sva[10]), .I4 (\z_out_2(10)  ), .I5 (nx28350z2)) ;
         defparam ix47647z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix47647z62756 (.O (nx47647z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[21]), .I4 (\z_out_2(10)  
         )) ;
         defparam ix47647z62756.INIT = 32'hFEEEF000;
    LUT6 ix28341z61890 (.O (nx28341z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[22]), .I3 (
         conv_core_inst_jj_sva[9]), .I4 (\z_out_2(9)  ), .I5 (nx28350z2)) ;
         defparam ix28341z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28341z62756 (.O (nx28341z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[22]), .I4 (\z_out_2(9)  )
         ) ;
         defparam ix28341z62756.INIT = 32'hFEEEF000;
    LUT6 ix28342z61890 (.O (nx28342z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[23]), .I3 (
         conv_core_inst_jj_sva[8]), .I4 (\z_out_2(8)  ), .I5 (nx28350z2)) ;
         defparam ix28342z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28342z62756 (.O (nx28342z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[23]), .I4 (\z_out_2(8)  )
         ) ;
         defparam ix28342z62756.INIT = 32'hFEEEF000;
    LUT6 ix28343z61890 (.O (nx28343z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[24]), .I3 (
         conv_core_inst_jj_sva[7]), .I4 (\z_out_2(7)  ), .I5 (nx28350z2)) ;
         defparam ix28343z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28343z62756 (.O (nx28343z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[24]), .I4 (\z_out_2(7)  )
         ) ;
         defparam ix28343z62756.INIT = 32'hFEEEF000;
    LUT6 ix28344z61890 (.O (nx28344z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[25]), .I3 (
         conv_core_inst_jj_sva[6]), .I4 (\z_out_2(6)  ), .I5 (nx28350z2)) ;
         defparam ix28344z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28344z62756 (.O (nx28344z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[25]), .I4 (\z_out_2(6)  )
         ) ;
         defparam ix28344z62756.INIT = 32'hFEEEF000;
    LUT6 ix28345z61890 (.O (nx28345z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[26]), .I3 (
         conv_core_inst_jj_sva[5]), .I4 (\z_out_2(5)  ), .I5 (nx28350z2)) ;
         defparam ix28345z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28345z62756 (.O (nx28345z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[26]), .I4 (\z_out_2(5)  )
         ) ;
         defparam ix28345z62756.INIT = 32'hFEEEF000;
    LUT6 ix28346z61890 (.O (nx28346z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[27]), .I3 (
         conv_core_inst_jj_sva[4]), .I4 (\z_out_2(4)  ), .I5 (nx28350z2)) ;
         defparam ix28346z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28346z62756 (.O (nx28346z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[27]), .I4 (\z_out_2(4)  )
         ) ;
         defparam ix28346z62756.INIT = 32'hFEEEF000;
    LUT6 ix28347z61890 (.O (nx28347z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[28]), .I3 (
         conv_core_inst_jj_sva[3]), .I4 (\z_out_2(3)  ), .I5 (nx28350z2)) ;
         defparam ix28347z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28347z62756 (.O (nx28347z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[28]), .I4 (\z_out_2(3)  )
         ) ;
         defparam ix28347z62756.INIT = 32'hFEEEF000;
    LUT6 ix28348z61890 (.O (nx28348z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[29]), .I3 (
         conv_core_inst_jj_sva[2]), .I4 (\z_out_2(2)  ), .I5 (nx28350z2)) ;
         defparam ix28348z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28348z62756 (.O (nx28348z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[29]), .I4 (\z_out_2(2)  )
         ) ;
         defparam ix28348z62756.INIT = 32'hFEEEF000;
    LUT6 ix28349z61890 (.O (nx28349z2), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[30]), .I3 (
         conv_core_inst_jj_sva[1]), .I4 (\z_out_2(1)  ), .I5 (nx28350z2)) ;
         defparam ix28349z61890.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28349z62756 (.O (nx28349z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[30]), .I4 (\z_out_2(1)  )
         ) ;
         defparam ix28349z62756.INIT = 32'hFEEEF000;
    LUT6 ix28350z61891 (.O (nx28350z1), .I0 (\fsm_output(5)  ), .I1 (
         \fsm_output(3)  ), .I2 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[31]), .I3 (
         conv_core_inst_jj_sva[0]), .I4 (\z_out_2(0)  ), .I5 (nx28350z2)) ;
         defparam ix28350z61891.INIT = 64'hECA0ECA0FFFFECA0;
    LUT5 ix28350z62758 (.O (nx28350z4), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(5)  ), .I3 (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[31]), .I4 (\z_out_2(0)  )
         ) ;
         defparam ix28350z62758.INIT = 32'hFEEEF000;
    LUT2 ix28350z1317 (.O (nx28350z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  )) ;
         defparam ix28350z1317.INIT = 4'h1;
    LUT3 ix39521z1427 (.O (nx39521z2), .I0 (\for_for_for_for_n_4_0_sva(4)  ), .I1 (
         nx39520z4), .I2 (nx39517z4)) ;
         defparam ix39521z1427.INIT = 8'h71;
    LUT6 ix39520z27325 (.O (nx39520z3), .I0 (\for_for_for_for_n_4_0_sva(4)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4]), .I2 (nx39517z1), .I3 (
         nx39520z4), .I4 (nx39519z4), .I5 (nx39517z4)) ;
         defparam ix39520z27325.INIT = 64'h59A69A65A659659A;
    LUT3 ix39520z1526 (.O (nx39520z2), .I0 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4]), .I1 (nx39517z1), .I2 (
         nx39519z4)) ;
         defparam ix39520z1526.INIT = 8'hD4;
    LUT5 ix39519z28600 (.O (nx39519z3), .I0 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4]), .I1 (
         \for_for_for_for_n_4_0_sva(2)  ), .I2 (nx39517z1), .I3 (nx39519z4), .I4 (
         nx39518z4)) ;
         defparam ix39519z28600.INIT = 32'hA9566A95;
    LUT3 ix39519z1526 (.O (nx39519z2), .I0 (\for_for_for_for_n_4_0_sva(2)  ), .I1 (
         nx39517z1), .I2 (nx39518z4)) ;
         defparam ix39519z1526.INIT = 8'hD4;
    LUT5 ix39518z28600 (.O (nx39518z3), .I0 (\for_for_for_for_n_4_0_sva(2)  ), .I1 (
         \for_for_for_for_n_4_0_sva(1)  ), .I2 (nx39517z1), .I3 (nx39518z4), .I4 (
         nx39517z6)) ;
         defparam ix39518z28600.INIT = 32'hA9566A95;
    LUT3 ix39518z1526 (.O (nx39518z2), .I0 (\for_for_for_for_n_4_0_sva(1)  ), .I1 (
         nx39517z1), .I2 (nx39517z6)) ;
         defparam ix39518z1526.INIT = 8'hD4;
    LUT6 ix39517z39882 (.O (nx39517z5), .I0 (\for_for_for_for_n_4_0_sva(1)  ), .I1 (
         \for_for_for_for_n_4_0_sva(0)  ), .I2 (nx39517z1), .I3 (nx39517z3), .I4 (
         nx39517z6), .I5 (nx39517z4)) ;
         defparam ix39517z39882.INIT = 64'hA5695A96695A96A5;
    LUT3 ix39517z1527 (.O (nx39517z2), .I0 (\for_for_for_for_n_4_0_sva(0)  ), .I1 (
         nx39517z3), .I2 (nx39517z4)) ;
         defparam ix39517z1527.INIT = 8'hD4;
    LUT4 ix50045z39820 (.O (nx50045z2), .I0 (nx39517z1), .I1 (nx39517z4), .I2 (
         \for_for_for_for_n_4_0_sva(0)  ), .I3 (nx39517z3)) ;
         defparam ix50045z39820.INIT = 16'h9669;
    LUT2 ix48536z1323 (.O (nx48536z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[30]), .I1 (
         conv_core_inst_rows_1_sva_2[1])) ;
         defparam ix48536z1323.INIT = 4'h9;
    LUT2 ix49524z1323 (.O (nx49524z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[29]), .I1 (
         conv_core_inst_rows_1_sva_2[2])) ;
         defparam ix49524z1323.INIT = 4'h9;
    LUT2 ix49525z1323 (.O (nx49525z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[28]), .I1 (
         conv_core_inst_rows_1_sva_2[3])) ;
         defparam ix49525z1323.INIT = 4'h9;
    LUT2 ix49526z1323 (.O (nx49526z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[27]), .I1 (
         conv_core_inst_rows_1_sva_2[4])) ;
         defparam ix49526z1323.INIT = 4'h9;
    LUT2 ix49527z1323 (.O (nx49527z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[26]), .I1 (
         conv_core_inst_rows_1_sva_2[5])) ;
         defparam ix49527z1323.INIT = 4'h9;
    LUT2 ix49528z1323 (.O (nx49528z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[25]), .I1 (
         conv_core_inst_rows_1_sva_2[6])) ;
         defparam ix49528z1323.INIT = 4'h9;
    LUT2 ix49529z1323 (.O (nx49529z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[24]), .I1 (
         conv_core_inst_rows_1_sva_2[7])) ;
         defparam ix49529z1323.INIT = 4'h9;
    LUT2 ix49530z1323 (.O (nx49530z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[23]), .I1 (
         conv_core_inst_rows_1_sva_2[8])) ;
         defparam ix49530z1323.INIT = 4'h9;
    LUT2 ix49531z1323 (.O (nx49531z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[22]), .I1 (
         conv_core_inst_rows_1_sva_2[9])) ;
         defparam ix49531z1323.INIT = 4'h9;
    LUT2 ix49532z1323 (.O (nx49532z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[21]), .I1 (
         conv_core_inst_rows_1_sva_2[10])) ;
         defparam ix49532z1323.INIT = 4'h9;
    LUT2 ix49533z1323 (.O (nx49533z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[20]), .I1 (
         conv_core_inst_rows_1_sva_2[11])) ;
         defparam ix49533z1323.INIT = 4'h9;
    LUT2 ix50521z1323 (.O (nx50521z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[19]), .I1 (
         conv_core_inst_rows_1_sva_2[12])) ;
         defparam ix50521z1323.INIT = 4'h9;
    LUT2 ix50522z1323 (.O (nx50522z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[18]), .I1 (
         conv_core_inst_rows_1_sva_2[13])) ;
         defparam ix50522z1323.INIT = 4'h9;
    LUT2 ix50523z1323 (.O (nx50523z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[17]), .I1 (
         conv_core_inst_rows_1_sva_2[14])) ;
         defparam ix50523z1323.INIT = 4'h9;
    LUT2 ix50524z1323 (.O (nx50524z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[16]), .I1 (
         conv_core_inst_rows_1_sva_2[15])) ;
         defparam ix50524z1323.INIT = 4'h9;
    LUT2 ix50525z1323 (.O (nx50525z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[15]), .I1 (
         conv_core_inst_rows_1_sva_2[16])) ;
         defparam ix50525z1323.INIT = 4'h9;
    LUT2 ix50526z1323 (.O (nx50526z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[14]), .I1 (
         conv_core_inst_rows_1_sva_2[17])) ;
         defparam ix50526z1323.INIT = 4'h9;
    LUT2 ix50527z1323 (.O (nx50527z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[13]), .I1 (
         conv_core_inst_rows_1_sva_2[18])) ;
         defparam ix50527z1323.INIT = 4'h9;
    LUT2 ix50528z1323 (.O (nx50528z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[12]), .I1 (
         conv_core_inst_rows_1_sva_2[19])) ;
         defparam ix50528z1323.INIT = 4'h9;
    LUT2 ix50529z1323 (.O (nx50529z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[11]), .I1 (
         conv_core_inst_rows_1_sva_2[20])) ;
         defparam ix50529z1323.INIT = 4'h9;
    LUT2 ix50530z1323 (.O (nx50530z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[10]), .I1 (
         conv_core_inst_rows_1_sva_2[21])) ;
         defparam ix50530z1323.INIT = 4'h9;
    LUT2 ix34270z1323 (.O (nx34270z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[9]), .I1 (
         conv_core_inst_rows_1_sva_2[22])) ;
         defparam ix34270z1323.INIT = 4'h9;
    LUT2 ix34269z1323 (.O (nx34269z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[8]), .I1 (
         conv_core_inst_rows_1_sva_2[23])) ;
         defparam ix34269z1323.INIT = 4'h9;
    LUT2 ix34268z1323 (.O (nx34268z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[7]), .I1 (
         conv_core_inst_rows_1_sva_2[24])) ;
         defparam ix34268z1323.INIT = 4'h9;
    LUT2 ix34267z1323 (.O (nx34267z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[6]), .I1 (
         conv_core_inst_rows_1_sva_2[25])) ;
         defparam ix34267z1323.INIT = 4'h9;
    LUT2 ix34266z1323 (.O (nx34266z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[5]), .I1 (
         conv_core_inst_rows_1_sva_2[26])) ;
         defparam ix34266z1323.INIT = 4'h9;
    LUT2 ix34265z1323 (.O (nx34265z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[4]), .I1 (
         conv_core_inst_rows_1_sva_2[27])) ;
         defparam ix34265z1323.INIT = 4'h9;
    LUT2 ix34264z1323 (.O (nx34264z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[3]), .I1 (
         conv_core_inst_rows_1_sva_2[28])) ;
         defparam ix34264z1323.INIT = 4'h9;
    LUT2 ix34263z1323 (.O (nx34263z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[2]), .I1 (
         conv_core_inst_rows_1_sva_2[29])) ;
         defparam ix34263z1323.INIT = 4'h9;
    LUT2 ix34262z1323 (.O (nx34262z2), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[1]), .I1 (
         conv_core_inst_rows_1_sva_2[30])) ;
         defparam ix34262z1323.INIT = 4'h9;
    LUT2 ix34261z1323 (.O (nx34261z1), .I0 (
         conv_core_inst_for_for_for_for_acc_3_tmp[0]), .I1 (
         conv_core_inst_rows_1_sva_2[31])) ;
         defparam ix34261z1323.INIT = 4'h9;
    (* HLUTNM = "LUT62_1_63" *)
    LUT3 ix7619z1483 (.O (nx7619z2), .I0 (conv_core_inst_for_i_sva[27]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix7619z1483.INIT = 8'hA9;
    LUT3 ix7618z1483 (.O (nx7618z2), .I0 (conv_core_inst_for_i_sva[26]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix7618z1483.INIT = 8'hA9;
    LUT3 ix6630z1483 (.O (nx6630z2), .I0 (conv_core_inst_for_i_sva[25]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6630z1483.INIT = 8'hA9;
    LUT3 ix6629z1483 (.O (nx6629z2), .I0 (conv_core_inst_for_i_sva[24]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6629z1483.INIT = 8'hA9;
    LUT3 ix6628z1483 (.O (nx6628z2), .I0 (conv_core_inst_for_i_sva[23]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6628z1483.INIT = 8'hA9;
    LUT3 ix6627z1483 (.O (nx6627z2), .I0 (conv_core_inst_for_i_sva[22]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6627z1483.INIT = 8'hA9;
    LUT3 ix6626z1483 (.O (nx6626z2), .I0 (conv_core_inst_for_i_sva[21]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6626z1483.INIT = 8'hA9;
    LUT3 ix6625z1483 (.O (nx6625z2), .I0 (conv_core_inst_for_i_sva[20]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6625z1483.INIT = 8'hA9;
    LUT3 ix6624z1483 (.O (nx6624z2), .I0 (conv_core_inst_for_i_sva[19]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6624z1483.INIT = 8'hA9;
    LUT3 ix6623z1483 (.O (nx6623z2), .I0 (conv_core_inst_for_i_sva[18]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6623z1483.INIT = 8'hA9;
    LUT3 ix6622z1483 (.O (nx6622z2), .I0 (conv_core_inst_for_i_sva[17]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6622z1483.INIT = 8'hA9;
    LUT3 ix6621z1483 (.O (nx6621z2), .I0 (conv_core_inst_for_i_sva[16]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix6621z1483.INIT = 8'hA9;
    LUT3 ix5633z1483 (.O (nx5633z2), .I0 (conv_core_inst_for_i_sva[15]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix5633z1483.INIT = 8'hA9;
    LUT3 ix5632z1483 (.O (nx5632z2), .I0 (conv_core_inst_for_i_sva[14]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix5632z1483.INIT = 8'hA9;
    LUT3 ix5631z1483 (.O (nx5631z2), .I0 (conv_core_inst_for_i_sva[13]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix5631z1483.INIT = 8'hA9;
    LUT3 ix5630z1483 (.O (nx5630z2), .I0 (conv_core_inst_for_i_sva[12]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix5630z1483.INIT = 8'hA9;
    LUT3 ix5629z1483 (.O (nx5629z2), .I0 (conv_core_inst_for_i_sva[11]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix5629z1483.INIT = 8'hA9;
    LUT3 ix5628z1483 (.O (nx5628z2), .I0 (conv_core_inst_for_i_sva[10]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix5628z1483.INIT = 8'hA9;
    LUT3 ix5627z1483 (.O (nx5627z2), .I0 (conv_core_inst_for_i_sva[9]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix5627z1483.INIT = 8'hA9;
    LUT3 ix5626z1483 (.O (nx5626z2), .I0 (conv_core_inst_for_i_sva[8]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix5626z1483.INIT = 8'hA9;
    LUT3 ix44834z1483 (.O (nx44834z2), .I0 (conv_core_inst_for_i_sva[7]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix44834z1483.INIT = 8'hA9;
    LUT3 ix44835z1483 (.O (nx44835z2), .I0 (conv_core_inst_for_i_sva[6]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix44835z1483.INIT = 8'hA9;
    LUT3 ix8911z1483 (.O (nx8911z2), .I0 (conv_core_inst_for_i_sva[5]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix8911z1483.INIT = 8'hA9;
    LUT3 ix8912z1483 (.O (nx8912z2), .I0 (conv_core_inst_for_i_sva[4]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix8912z1483.INIT = 8'hA9;
    LUT3 ix8913z1483 (.O (nx8913z2), .I0 (conv_core_inst_for_i_sva[3]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix8913z1483.INIT = 8'hA9;
    LUT3 ix8914z1483 (.O (nx8914z2), .I0 (conv_core_inst_for_i_sva[2]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix8914z1483.INIT = 8'hA9;
    LUT3 ix8915z1483 (.O (nx8915z2), .I0 (conv_core_inst_for_i_sva[1]), .I1 (
         nx20393z3), .I2 (nx18544z2)) ;
         defparam ix8915z1483.INIT = 8'hA9;
    LUT2 ix8917z1324 (.O (nx8917z2), .I0 (conv_core_inst_for_i_sva[28]), .I1 (
         nx18544z2)) ;
         defparam ix8917z1324.INIT = 4'h9;
    LUT2 ix63169z1323 (.O (nx63169z2), .I0 (\for_for_j_sva(3)  ), .I1 (
         conv_core_inst_for_for_for_for_n_4_0_sva[4])) ;
         defparam ix63169z1323.INIT = 4'h9;
    LUT4 ix6185z22323 (.O (nx6185z31), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[31]), .I3 (
         conv_core_inst_for_i_sva[31])) ;
         defparam ix6185z22323.INIT = 16'h51F3;
    LUT4 ix6185z22322 (.O (nx6185z30), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[30]), .I3 (
         conv_core_inst_for_i_sva[30])) ;
         defparam ix6185z22322.INIT = 16'h51F3;
    LUT4 ix6185z22321 (.O (nx6185z29), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[29]), .I3 (
         conv_core_inst_for_i_sva[29])) ;
         defparam ix6185z22321.INIT = 16'h51F3;
    LUT4 ix6185z22320 (.O (nx6185z28), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[28]), .I3 (
         \for_for_j_sva(3)  )) ;
         defparam ix6185z22320.INIT = 16'h51F3;
    LUT4 ix6185z22319 (.O (nx6185z27), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[27]), .I3 (
         \for_for_j_sva(4)  )) ;
         defparam ix6185z22319.INIT = 16'h51F3;
    LUT4 ix6185z22318 (.O (nx6185z26), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[26]), .I3 (
         \for_for_j_sva(5)  )) ;
         defparam ix6185z22318.INIT = 16'h51F3;
    LUT4 ix6185z22317 (.O (nx6185z25), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[25]), .I3 (
         \for_for_j_sva(6)  )) ;
         defparam ix6185z22317.INIT = 16'h51F3;
    LUT4 ix6185z22316 (.O (nx6185z24), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[24]), .I3 (
         \for_for_j_sva(7)  )) ;
         defparam ix6185z22316.INIT = 16'h51F3;
    LUT4 ix6185z22315 (.O (nx6185z23), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[23]), .I3 (
         \for_for_j_sva(8)  )) ;
         defparam ix6185z22315.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_37" *)
    LUT4 ix6185z22314 (.O (nx6185z22), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[22]), .I3 (
         \for_for_j_sva(9)  )) ;
         defparam ix6185z22314.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_36" *)
    LUT4 ix6185z22313 (.O (nx6185z21), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[21]), .I3 (
         \for_for_j_sva(10)  )) ;
         defparam ix6185z22313.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_35" *)
    LUT4 ix6185z22312 (.O (nx6185z20), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[20]), .I3 (
         \for_for_j_sva(11)  )) ;
         defparam ix6185z22312.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_34" *)
    LUT4 ix6185z22311 (.O (nx6185z19), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[19]), .I3 (
         \for_for_j_sva(12)  )) ;
         defparam ix6185z22311.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_33" *)
    LUT4 ix6185z22310 (.O (nx6185z18), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[18]), .I3 (
         \for_for_j_sva(13)  )) ;
         defparam ix6185z22310.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_32" *)
    LUT4 ix6185z22309 (.O (nx6185z17), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[17]), .I3 (
         \for_for_j_sva(14)  )) ;
         defparam ix6185z22309.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_31" *)
    LUT4 ix6185z22308 (.O (nx6185z16), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[16]), .I3 (
         \for_for_j_sva(15)  )) ;
         defparam ix6185z22308.INIT = 16'h51F3;
    LUT4 ix6185z22307 (.O (nx6185z15), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[15]), .I3 (
         \for_for_j_sva(16)  )) ;
         defparam ix6185z22307.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_30" *)
    LUT4 ix6185z22306 (.O (nx6185z14), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[14]), .I3 (
         \for_for_j_sva(17)  )) ;
         defparam ix6185z22306.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_29" *)
    LUT4 ix6185z22305 (.O (nx6185z13), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[13]), .I3 (
         \for_for_j_sva(18)  )) ;
         defparam ix6185z22305.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_28" *)
    LUT4 ix6185z22304 (.O (nx6185z12), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[12]), .I3 (
         \for_for_j_sva(19)  )) ;
         defparam ix6185z22304.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_27" *)
    LUT4 ix6185z22303 (.O (nx6185z11), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[11]), .I3 (
         \for_for_j_sva(20)  )) ;
         defparam ix6185z22303.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_26" *)
    LUT4 ix6185z22302 (.O (nx6185z10), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[10]), .I3 (
         \for_for_j_sva(21)  )) ;
         defparam ix6185z22302.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_25" *)
    LUT4 ix6185z22301 (.O (nx6185z9), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[9]), .I3 (
         \for_for_j_sva(22)  )) ;
         defparam ix6185z22301.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_24" *)
    LUT4 ix6185z22300 (.O (nx6185z8), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[8]), .I3 (
         \for_for_j_sva(23)  )) ;
         defparam ix6185z22300.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_23" *)
    LUT4 ix6185z22299 (.O (nx6185z7), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[7]), .I3 (
         \for_for_j_sva(24)  )) ;
         defparam ix6185z22299.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_22" *)
    LUT4 ix6185z22298 (.O (nx6185z6), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[6]), .I3 (
         \for_for_j_sva(25)  )) ;
         defparam ix6185z22298.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_21" *)
    LUT4 ix6185z22297 (.O (nx6185z5), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[5]), .I3 (
         \for_for_j_sva(26)  )) ;
         defparam ix6185z22297.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_20" *)
    LUT4 ix6185z22296 (.O (nx6185z4), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[4]), .I3 (
         \for_for_j_sva(27)  )) ;
         defparam ix6185z22296.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_19" *)
    LUT4 ix6185z22295 (.O (nx6185z3), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[3]), .I3 (
         \for_for_j_sva(28)  )) ;
         defparam ix6185z22295.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_18" *)
    LUT4 ix6185z22294 (.O (nx6185z2), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[2]), .I3 (
         \for_for_j_sva(29)  )) ;
         defparam ix6185z22294.INIT = 16'h51F3;
    (* HLUTNM = "LUT62_1_4" *)
    LUT4 ix6185z22293 (.O (nx6185z1), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(1)  ), .I2 (conv_core_inst_cols_1_sva_1[1]), .I3 (
         \for_for_j_sva(30)  )) ;
         defparam ix6185z22293.INIT = 16'h51F3;
    LUT2 ix23435z1321 (.O (px1534), .I0 (\fsm_output(4)  ), .I1 (
         for_for_for_for_if_for_for_for_for_if_and_2_itm)) ;
         defparam ix23435z1321.INIT = 4'h7;
    (* HLUTNM = "LUT62_1_45" *)
    LUT3 ix23434z1530 (.O (px1535), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[0]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[13])) ;
         defparam ix23434z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_45" *)
    LUT3 ix23433z1530 (.O (px1536), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[1]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[12])) ;
         defparam ix23433z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_44" *)
    LUT3 ix23432z1530 (.O (px1537), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[2]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[11])) ;
         defparam ix23432z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_44" *)
    LUT3 ix23431z1530 (.O (px1538), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[3]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[10])) ;
         defparam ix23431z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_43" *)
    LUT3 ix23430z1530 (.O (px1539), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[4]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[9])) ;
         defparam ix23430z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_43" *)
    LUT3 ix22442z1530 (.O (px1540), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[5]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[8])) ;
         defparam ix22442z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_42" *)
    LUT3 ix22441z1530 (.O (px1541), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[6]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[7])) ;
         defparam ix22441z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_42" *)
    LUT3 ix22440z1530 (.O (px1542), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[7]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[6])) ;
         defparam ix22440z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_41" *)
    LUT3 ix22439z1530 (.O (px1543), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[8]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[5])) ;
         defparam ix22439z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_41" *)
    LUT3 ix22438z1530 (.O (px1544), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[9]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[4])) ;
         defparam ix22438z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_40" *)
    LUT3 ix22437z1530 (.O (px1545), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[10]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[3])) ;
         defparam ix22437z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_40" *)
    LUT3 ix22436z1530 (.O (px1546), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[11]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[2])) ;
         defparam ix22436z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_39" *)
    LUT3 ix22435z1530 (.O (px1547), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[12]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[1])) ;
         defparam ix22435z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_39" *)
    LUT3 ix22434z1530 (.O (px1548), .I0 (\fsm_output(5)  ), .I1 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva_1[13]), .I2 (
         conv_core_inst_for_for_for_for_if_acc_psp_sva[0])) ;
         defparam ix22434z1530.INIT = 8'hD8;
    LUT6 ix22433z1313 (.O (px1549), .I0 (\fsm_output(3)  ), .I1 (
         conv_core_inst_for_for_for_for_acc_3_tmp[31]), .I2 (
         conv_core_inst_rows_1_sva_2[0]), .I3 (conv_core_inst_jj_sva[31]), .I4 (
         \z_out_1(32)  ), .I5 (nx60570z2)) ;
         defparam ix22433z1313.INIT = 64'hFFFFFFFFFFFDFFFF;
    (* HLUTNM = "LUT62_1_9" *)
    LUT2 ix21445z1321 (.O (px1550), .I0 (\fsm_output(5)  ), .I1 (
         for_for_for_for_if_for_for_for_for_if_and_2_itm)) ;
         defparam ix21445z1321.INIT = 4'h7;
    LUT5 ix49642z54064 (.O (nx49642z6), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(5)  ), .I2 (conv_core_inst_cols_1_sva_1[0]), .I3 (
         \z_out_4(31)  ), .I4 (\fsm_output(3)  )) ;
         defparam ix49642z54064.INIT = 32'hCF0FCE0A;
    DSP48E1 z_out_4_multu32_0_p_mult0_DSP48E1_0 (.BCOUT ({nx18281z16,nx18281z17,
            nx18281z18,nx18281z19,nx18281z20,nx18281z21,nx18281z22,nx18281z23,
            nx18281z24,nx18281z25,nx18281z26,nx18281z27,nx18281z28,nx18281z29,
            nx18281z30,nx18281z31,nx18281z32,nx18281z33}), .P ({\$dummy [0],
            \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
            \$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],\$dummy [10],
            \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],\$dummy [15],
            \$dummy [16],\$dummy [17],\$dummy [18],\$dummy [19],\$dummy [20],
            \$dummy [21],\$dummy [22],\$dummy [23],\$dummy [24],\$dummy [25],
            \$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29],\$dummy [30],
            \z_out_4(16)  ,\z_out_4(15)  ,\z_out_4(14)  ,\z_out_4(13)  ,
            \z_out_4(12)  ,\z_out_4(11)  ,\z_out_4(10)  ,\z_out_4(9)  ,
            \z_out_4(8)  ,\z_out_4(7)  ,\z_out_4(6)  ,\z_out_4(5)  ,\z_out_4(4)  
            ,\z_out_4(3)  ,\z_out_4(2)  ,\z_out_4(1)  ,\z_out_4(0)  }), .PCOUT (
            {nx18281z34,nx18281z35,nx18281z36,nx18281z37,nx18281z38,nx18281z39,
            nx18281z40,nx18281z41,nx18281z42,nx18281z43,nx18281z44,nx18281z45,
            nx18281z46,nx18281z47,nx18281z48,nx18281z49,nx18281z50,nx18281z51,
            nx18281z52,nx18281z53,nx18281z54,nx18281z55,nx18281z56,nx18281z57,
            nx18281z58,nx18281z59,nx18281z60,nx18281z61,nx18281z62,nx18281z63,
            nx18281z64,nx18281z65,nx18281z66,nx18281z67,nx18281z68,nx18281z69,
            nx18281z70,nx18281z71,nx18281z72,nx18281z73,nx18281z74,nx18281z75,
            nx18281z76,nx18281z77,nx18281z78,nx18281z79,nx18281z80,nx18281z81})
            , .A ({px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,nx30685z1,nx30685z2,nx30685z3,
            nx30685z4,nx30685z5,nx30685z6,nx30685z7,nx30685z8,nx30685z9,
            nx30685z10,nx30685z11,nx30685z12,nx30685z13,nx30685z14,nx30685z15,
            nx30685z16,nx30685z17}), .ALUMODE ({px1140,px1140,px1140,px1140}), .B (
            {px1140,nx30685z18,nx30685z19,nx30685z20,nx30685z21,nx30685z22,
            nx30685z23,nx30685z24,nx30685z25,nx30685z26,nx30685z27,nx30685z28,
            nx30685z29,nx30685z30,nx30685z31,nx30685z32,nx30685z33,nx30685z34})
            , .C ({px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140}), .CARRYCASCIN (px1140), .CARRYIN (
            px1140), .CARRYINSEL ({px1140,px1140,px1140}), .CEA1 (px1140), .CEA2 (
            px1140), .CEAD (px1140), .CEALUMODE (px1140), .CEB1 (px1140), .CEB2 (
            px1140), .CEC (px1140), .CECARRYIN (px1140), .CECTRL (px1140), .CED (
            px1140), .CEINMODE (px1140), .CEM (px1140), .CEP (px1140), .CLK (
            px1140), .D ({px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140}), .INMODE (
            {px1140,px1140,px1140,px1140,px1140}), .MULTSIGNIN (px1551), .OPMODE (
            {px1140,px1140,px1140,px1140,px1551,px1140,px1551}), .RSTA (px1140)
            , .RSTALLCARRYIN (px1140), .RSTALUMODE (px1140), .RSTB (px1140), .RSTC (
            px1140), .RSTCTRL (px1140), .RSTD (px1140), .RSTINMODE (px1140), .RSTM (
            px1140), .RSTP (px1140)) ;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.ACASCREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.ADREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.ALUMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.AREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.AUTORESET_PATDET = "NO_RESET";
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.A_INPUT = "DIRECT";
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.BCASCREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.BREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.B_INPUT = "DIRECT";
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.CARRYINREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.CARRYINSELREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.CREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.DREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.INMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.MREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.OPMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.PREG = 0;
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.SEL_MASK = "MASK";
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.SEL_PATTERN = "PATTERN";
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.USE_DPORT = "FALSE";
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.USE_MULT = "MULTIPLY";
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.USE_PATTERN_DETECT = "NO_PATDET";
            defparam z_out_4_multu32_0_p_mult0_DSP48E1_0.USE_SIMD = "ONE48";
    DSP48E1 z_out_4_multu32_0_p_mult1_DSP48E1_1 (.PCOUT ({nx63825z16,nx63825z17,
            nx63825z18,nx63825z19,nx63825z20,nx63825z21,nx63825z22,nx63825z23,
            nx63825z24,nx63825z25,nx63825z26,nx63825z27,nx63825z28,nx63825z29,
            nx63825z30,nx63825z31,nx63825z32,nx63825z33,nx63825z34,nx63825z35,
            nx63825z36,nx63825z37,nx63825z38,nx63825z39,nx63825z40,nx63825z41,
            nx63825z42,nx63825z43,nx63825z44,nx63825z45,nx63825z46,nx63825z47,
            nx63825z48,nx63825z49,nx63825z50,nx63825z51,nx63825z52,nx63825z53,
            nx63825z54,nx63825z55,nx63825z56,nx63825z57,nx63825z58,nx63825z59,
            nx63825z60,nx63825z61,nx63825z62,nx63825z63}), .A ({px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,nx18281z1,nx18281z2,nx18281z3,nx18281z4,
            nx18281z5,nx18281z6,nx18281z7,nx18281z8,nx18281z9,nx18281z10,
            nx18281z11,nx18281z12,nx18281z13,nx18281z14,nx18281z15}), .ALUMODE (
            {px1140,px1140,px1140,px1140}), .BCIN ({nx18281z16,nx18281z17,
            nx18281z18,nx18281z19,nx18281z20,nx18281z21,nx18281z22,nx18281z23,
            nx18281z24,nx18281z25,nx18281z26,nx18281z27,nx18281z28,nx18281z29,
            nx18281z30,nx18281z31,nx18281z32,nx18281z33}), .C ({px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140}), .CARRYCASCIN (px1140), .CARRYIN (px1140), .CARRYINSEL ({
            px1140,px1140,px1140}), .CEA1 (px1140), .CEA2 (px1140), .CEAD (
            px1140), .CEALUMODE (px1140), .CEB1 (px1140), .CEB2 (px1140), .CEC (
            px1140), .CECARRYIN (px1140), .CECTRL (px1140), .CED (px1140), .CEINMODE (
            px1140), .CEM (px1140), .CEP (px1140), .CLK (px1140), .D ({px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140}), .INMODE ({px1140,px1140
            ,px1140,px1140,px1140}), .MULTSIGNIN (px1551), .OPMODE ({px1551,
            px1140,px1551,px1140,px1551,px1140,px1551}), .PCIN ({nx18281z34,
            nx18281z35,nx18281z36,nx18281z37,nx18281z38,nx18281z39,nx18281z40,
            nx18281z41,nx18281z42,nx18281z43,nx18281z44,nx18281z45,nx18281z46,
            nx18281z47,nx18281z48,nx18281z49,nx18281z50,nx18281z51,nx18281z52,
            nx18281z53,nx18281z54,nx18281z55,nx18281z56,nx18281z57,nx18281z58,
            nx18281z59,nx18281z60,nx18281z61,nx18281z62,nx18281z63,nx18281z64,
            nx18281z65,nx18281z66,nx18281z67,nx18281z68,nx18281z69,nx18281z70,
            nx18281z71,nx18281z72,nx18281z73,nx18281z74,nx18281z75,nx18281z76,
            nx18281z77,nx18281z78,nx18281z79,nx18281z80,nx18281z81}), .RSTA (
            px1140), .RSTALLCARRYIN (px1140), .RSTALUMODE (px1140), .RSTB (
            px1140), .RSTC (px1140), .RSTCTRL (px1140), .RSTD (px1140), .RSTINMODE (
            px1140), .RSTM (px1140), .RSTP (px1140)) ;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.ACASCREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.ADREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.ALUMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.AREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.AUTORESET_PATDET = "NO_RESET";
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.A_INPUT = "DIRECT";
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.BCASCREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.BREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.B_INPUT = "CASCADE";
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.CARRYINREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.CARRYINSELREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.CREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.DREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.INMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.MREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.OPMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.PREG = 0;
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.SEL_MASK = "MASK";
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.SEL_PATTERN = "PATTERN";
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.USE_DPORT = "FALSE";
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.USE_MULT = "MULTIPLY";
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.USE_PATTERN_DETECT = "NO_PATDET";
            defparam z_out_4_multu32_0_p_mult1_DSP48E1_1.USE_SIMD = "ONE48";
    DSP48E1 z_out_4_multu32_0_p_mult2_DSP48E1_2 (.P ({\$dummy [31],\$dummy [32],
            \$dummy [33],\$dummy [34],\$dummy [35],\$dummy [36],\$dummy [37],
            \$dummy [38],\$dummy [39],\$dummy [40],\$dummy [41],\$dummy [42],
            \$dummy [43],\$dummy [44],\$dummy [45],\$dummy [46],\$dummy [47],
            \$dummy [48],\$dummy [49],\$dummy [50],\$dummy [51],\$dummy [52],
            \$dummy [53],\$dummy [54],\$dummy [55],\$dummy [56],\$dummy [57],
            \$dummy [58],\$dummy [59],\$dummy [60],\$dummy [61],\$dummy [62],
            \$dummy [63],\z_out_4(31)  ,\z_out_4(30)  ,\z_out_4(29)  ,
            \z_out_4(28)  ,\z_out_4(27)  ,\z_out_4(26)  ,\z_out_4(25)  ,
            \z_out_4(24)  ,\z_out_4(23)  ,\z_out_4(22)  ,\z_out_4(21)  ,
            \z_out_4(20)  ,\z_out_4(19)  ,\z_out_4(18)  ,
            conv_core_inst_z_out_4[31]}), .A ({px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            nx30685z1,nx30685z2,nx30685z3,nx30685z4,nx30685z5,nx30685z6,
            nx30685z7,nx30685z8,nx30685z9,nx30685z10,nx30685z11,nx30685z12,
            nx30685z13,nx30685z14,nx30685z15,nx30685z16,nx30685z17}), .ALUMODE (
            {px1140,px1140,px1140,px1140}), .B ({px1140,px1140,px1140,nx63825z1,
            nx63825z2,nx63825z3,nx63825z4,nx63825z5,nx63825z6,nx63825z7,
            nx63825z8,nx63825z9,nx63825z10,nx63825z11,nx63825z12,nx63825z13,
            nx63825z14,nx63825z15}), .C ({px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140}), .CARRYCASCIN (
            px1140), .CARRYIN (px1140), .CARRYINSEL ({px1140,px1140,px1140}), .CEA1 (
            px1140), .CEA2 (px1140), .CEAD (px1140), .CEALUMODE (px1140), .CEB1 (
            px1140), .CEB2 (px1140), .CEC (px1140), .CECARRYIN (px1140), .CECTRL (
            px1140), .CED (px1140), .CEINMODE (px1140), .CEM (px1140), .CEP (
            px1140), .CLK (px1140), .D ({px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,px1140,
            px1140,px1140}), .INMODE ({px1140,px1140,px1140,px1140,px1140}), .MULTSIGNIN (
            px1551), .OPMODE ({px1140,px1140,px1551,px1140,px1551,px1140,px1551}
            ), .PCIN ({nx63825z16,nx63825z17,nx63825z18,nx63825z19,nx63825z20,
            nx63825z21,nx63825z22,nx63825z23,nx63825z24,nx63825z25,nx63825z26,
            nx63825z27,nx63825z28,nx63825z29,nx63825z30,nx63825z31,nx63825z32,
            nx63825z33,nx63825z34,nx63825z35,nx63825z36,nx63825z37,nx63825z38,
            nx63825z39,nx63825z40,nx63825z41,nx63825z42,nx63825z43,nx63825z44,
            nx63825z45,nx63825z46,nx63825z47,nx63825z48,nx63825z49,nx63825z50,
            nx63825z51,nx63825z52,nx63825z53,nx63825z54,nx63825z55,nx63825z56,
            nx63825z57,nx63825z58,nx63825z59,nx63825z60,nx63825z61,nx63825z62,
            nx63825z63}), .RSTA (px1140), .RSTALLCARRYIN (px1140), .RSTALUMODE (
            px1140), .RSTB (px1140), .RSTC (px1140), .RSTCTRL (px1140), .RSTD (
            px1140), .RSTINMODE (px1140), .RSTM (px1140), .RSTP (px1140)) ;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.ACASCREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.ADREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.ALUMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.AREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.AUTORESET_PATDET = "NO_RESET";
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.A_INPUT = "DIRECT";
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.BCASCREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.BREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.B_INPUT = "DIRECT";
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.CARRYINREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.CARRYINSELREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.CREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.DREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.INMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.MREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.OPMODEREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.PREG = 0;
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.SEL_MASK = "MASK";
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.SEL_PATTERN = "PATTERN";
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.USE_DPORT = "FALSE";
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.USE_MULT = "MULTIPLY";
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.USE_PATTERN_DETECT = "NO_PATDET";
            defparam z_out_4_multu32_0_p_mult2_DSP48E1_2.USE_SIMD = "ONE48";
    LUT6 ix14411z44834 (.O (nx14411z1), .I0 (nx12614z1), .I1 (nx14411z2), .I2 (
         \z_out_1(32)  ), .I3 (\fsm_output(7)  ), .I4 (\fsm_output(1)  ), .I5 (
         \fsm_output(8)  )) ;
         defparam ix14411z44834.INIT = 64'hFAF0FAF0EECCAA00;
    LUT6 ix21390z1314 (.O (nx21390z1), .I0 (nx13414z2), .I1 (nx22387z2), .I2 (
         nx21390z2), .I3 (\z_out_1(32)  ), .I4 (\fsm_output(1)  ), .I5 (
         \fsm_output(8)  )) ;
         defparam ix21390z1314.INIT = 64'h00FF00FFF8F80000;
    LUT6 ix22387z1314 (.O (nx22387z1), .I0 (nx13414z2), .I1 (nx22387z2), .I2 (
         nx21390z2), .I3 (\z_out_1(32)  ), .I4 (\fsm_output(0)  ), .I5 (
         \fsm_output(9)  )) ;
         defparam ix22387z1314.INIT = 64'h00FF00FFF8F80000;
    LUT6 ix13414z1314 (.O (nx13414z1), .I0 (nx13414z2), .I1 (nx22387z2), .I2 (
         nx21390z2), .I3 (\z_out_1(32)  ), .I4 (\fsm_output(0)  ), .I5 (
         \fsm_output(9)  )) ;
         defparam ix13414z1314.INIT = 64'hFF00FF0007070000;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_0 (.O (nx23676z1), .CI (
          px1140), .DI (\z_out_4(0)  ), .S (nx23677z1)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_1 (.O (nx23675z1), .CI (
          nx23676z1), .DI (\z_out_4(1)  ), .S (nx23676z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_2 (.O (nx23674z1), .CI (
          nx23675z1), .DI (\z_out_4(2)  ), .S (nx23675z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_3 (.O (nx23673z1), .CI (
          nx23674z1), .DI (\z_out_4(3)  ), .S (nx23674z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_4 (.O (nx23672z1), .CI (
          nx23673z1), .DI (\z_out_4(4)  ), .S (nx23673z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_5 (.O (nx23671z1), .CI (
          nx23672z1), .DI (\z_out_4(5)  ), .S (nx23672z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_6 (.O (nx23670z1), .CI (
          nx23671z1), .DI (\z_out_4(6)  ), .S (nx23671z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_7 (.O (nx23669z1), .CI (
          nx23670z1), .DI (\z_out_4(7)  ), .S (nx23670z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_8 (.O (nx23668z1), .CI (
          nx23669z1), .DI (\z_out_4(8)  ), .S (nx23669z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_9 (.O (nx11964z1), .CI (
          nx23668z1), .DI (\z_out_4(9)  ), .S (nx23668z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_10 (.O (nx11963z1), .CI (
          nx11964z1), .DI (\z_out_4(10)  ), .S (nx11964z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_11 (.O (nx11962z1), .CI (
          nx11963z1), .DI (\z_out_4(11)  ), .S (nx11963z2)) ;
    MUXCY for_for_for_for_if_acc_psp_sva_add14_0_muxcy_12 (.O (nx11961z1), .CI (
          nx11962z1), .DI (\z_out_4(12)  ), .S (nx11962z2)) ;
    MUXCY jj_sva_add32_2_muxcy_0 (.O (nx63167z1), .CI (px1140), .DI (
          \for_for_for_for_n_4_0_sva(0)  ), .S (nx63166z2)) ;
    MUXCY jj_sva_add32_2_muxcy_1 (.O (nx63168z1), .CI (nx63167z1), .DI (
          \for_for_for_for_n_4_0_sva(1)  ), .S (nx63167z2)) ;
    MUXCY jj_sva_add32_2_muxcy_2 (.O (nx63169z1), .CI (nx63168z1), .DI (
          \for_for_for_for_n_4_0_sva(2)  ), .S (nx63168z2)) ;
    MUXCY jj_sva_add32_2_muxcy_3 (.O (nx63170z1), .CI (nx63169z1), .DI (
          \kernel_rsci_addr_d_0n0s2(3)  ), .S (nx63169z2)) ;
    MUXCY jj_sva_add32_2_muxcy_4 (.O (nx63171z1), .CI (nx63170z1), .DI (
          \for_for_j_sva(4)  ), .S (nx63170z2)) ;
    MUXCY jj_sva_add32_2_muxcy_5 (.O (nx63172z1), .CI (nx63171z1), .DI (
          \for_for_j_sva(5)  ), .S (nx63171z2)) ;
    MUXCY jj_sva_add32_2_muxcy_6 (.O (nx63173z1), .CI (nx63172z1), .DI (
          \for_for_j_sva(6)  ), .S (nx63172z2)) ;
    MUXCY jj_sva_add32_2_muxcy_7 (.O (nx63174z1), .CI (nx63173z1), .DI (
          \for_for_j_sva(7)  ), .S (nx63173z2)) ;
    MUXCY jj_sva_add32_2_muxcy_8 (.O (nx63175z1), .CI (nx63174z1), .DI (
          \for_for_j_sva(8)  ), .S (nx63174z2)) ;
    MUXCY jj_sva_add32_2_muxcy_9 (.O (nx62987z1), .CI (nx63175z1), .DI (
          \for_for_j_sva(9)  ), .S (nx63175z2)) ;
    MUXCY jj_sva_add32_2_muxcy_10 (.O (nx62988z1), .CI (nx62987z1), .DI (
          \for_for_j_sva(10)  ), .S (nx62987z2)) ;
    MUXCY jj_sva_add32_2_muxcy_11 (.O (nx62989z1), .CI (nx62988z1), .DI (
          \for_for_j_sva(11)  ), .S (nx62988z2)) ;
    MUXCY jj_sva_add32_2_muxcy_12 (.O (nx62990z1), .CI (nx62989z1), .DI (
          \for_for_j_sva(12)  ), .S (nx62989z2)) ;
    MUXCY jj_sva_add32_2_muxcy_13 (.O (nx62991z1), .CI (nx62990z1), .DI (
          \for_for_j_sva(13)  ), .S (nx62990z2)) ;
    MUXCY jj_sva_add32_2_muxcy_14 (.O (nx62992z1), .CI (nx62991z1), .DI (
          \for_for_j_sva(14)  ), .S (nx62991z2)) ;
    MUXCY jj_sva_add32_2_muxcy_15 (.O (nx62993z1), .CI (nx62992z1), .DI (
          \for_for_j_sva(15)  ), .S (nx62992z2)) ;
    MUXCY jj_sva_add32_2_muxcy_16 (.O (nx62994z1), .CI (nx62993z1), .DI (
          \for_for_j_sva(16)  ), .S (nx62993z2)) ;
    MUXCY jj_sva_add32_2_muxcy_17 (.O (nx62995z1), .CI (nx62994z1), .DI (
          \for_for_j_sva(17)  ), .S (nx62994z2)) ;
    MUXCY jj_sva_add32_2_muxcy_18 (.O (nx62996z1), .CI (nx62995z1), .DI (
          \for_for_j_sva(18)  ), .S (nx62995z2)) ;
    MUXCY jj_sva_add32_2_muxcy_19 (.O (nx63984z1), .CI (nx62996z1), .DI (
          \for_for_j_sva(19)  ), .S (nx62996z2)) ;
    MUXCY jj_sva_add32_2_muxcy_20 (.O (nx63985z1), .CI (nx63984z1), .DI (
          \for_for_j_sva(20)  ), .S (nx63984z2)) ;
    MUXCY jj_sva_add32_2_muxcy_21 (.O (nx63986z1), .CI (nx63985z1), .DI (
          \for_for_j_sva(21)  ), .S (nx63985z2)) ;
    MUXCY jj_sva_add32_2_muxcy_22 (.O (nx63987z1), .CI (nx63986z1), .DI (
          \for_for_j_sva(22)  ), .S (nx63986z2)) ;
    MUXCY jj_sva_add32_2_muxcy_23 (.O (nx63988z1), .CI (nx63987z1), .DI (
          \for_for_j_sva(23)  ), .S (nx63987z2)) ;
    MUXCY jj_sva_add32_2_muxcy_24 (.O (nx63989z1), .CI (nx63988z1), .DI (
          \for_for_j_sva(24)  ), .S (nx63988z2)) ;
    MUXCY jj_sva_add32_2_muxcy_25 (.O (nx63990z1), .CI (nx63989z1), .DI (
          \for_for_j_sva(25)  ), .S (nx63989z2)) ;
    MUXCY jj_sva_add32_2_muxcy_26 (.O (nx63991z1), .CI (nx63990z1), .DI (
          \for_for_j_sva(26)  ), .S (nx63990z2)) ;
    MUXCY jj_sva_add32_2_muxcy_27 (.O (nx63992z1), .CI (nx63991z1), .DI (
          \for_for_j_sva(27)  ), .S (nx63991z2)) ;
    MUXCY jj_sva_add32_2_muxcy_28 (.O (nx63993z1), .CI (nx63992z1), .DI (
          \for_for_j_sva(28)  ), .S (nx63992z2)) ;
    MUXCY jj_sva_add32_2_muxcy_29 (.O (nx64981z1), .CI (nx63993z1), .DI (
          \for_for_j_sva(29)  ), .S (nx63993z2)) ;
    MUXCY jj_sva_add32_2_muxcy_30 (.O (nx64982z1), .CI (nx64981z1), .DI (
          \for_for_j_sva(30)  ), .S (nx64981z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_0 (.O (nx8919z1), .CI (px1140)
          , .DI (nx12614z3), .S (nx8920z1)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_1 (.O (nx8918z1), .CI (
          nx8919z1), .DI (nx20538z2), .S (nx8919z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_2 (.O (nx8917z1), .CI (
          nx8918z1), .DI (nx19541z2), .S (nx8918z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_3 (.O (nx8916z1), .CI (
          nx8917z1), .DI (\for_for_for_acc_1_psp_sva_11n1s2(3)  ), .S (nx8917z2)
          ) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_4 (.O (nx8915z1), .CI (
          nx8916z1), .DI (conv_core_inst_for_i_sva[0]), .S (nx8916z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_5 (.O (nx8914z1), .CI (
          nx8915z1), .DI (conv_core_inst_for_i_sva[1]), .S (nx8915z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_6 (.O (nx8913z1), .CI (
          nx8914z1), .DI (conv_core_inst_for_i_sva[2]), .S (nx8914z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_7 (.O (nx8912z1), .CI (
          nx8913z1), .DI (conv_core_inst_for_i_sva[3]), .S (nx8913z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_8 (.O (nx8911z1), .CI (
          nx8912z1), .DI (conv_core_inst_for_i_sva[4]), .S (nx8912z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_9 (.O (nx44835z1), .CI (
          nx8911z1), .DI (conv_core_inst_for_i_sva[5]), .S (nx8911z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_10 (.O (nx44834z1), .CI (
          nx44835z1), .DI (conv_core_inst_for_i_sva[6]), .S (nx44835z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_11 (.O (nx5626z1), .CI (
          nx44834z1), .DI (conv_core_inst_for_i_sva[7]), .S (nx44834z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_12 (.O (nx5627z1), .CI (
          nx5626z1), .DI (conv_core_inst_for_i_sva[8]), .S (nx5626z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_13 (.O (nx5628z1), .CI (
          nx5627z1), .DI (conv_core_inst_for_i_sva[9]), .S (nx5627z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_14 (.O (nx5629z1), .CI (
          nx5628z1), .DI (conv_core_inst_for_i_sva[10]), .S (nx5628z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_15 (.O (nx5630z1), .CI (
          nx5629z1), .DI (conv_core_inst_for_i_sva[11]), .S (nx5629z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_16 (.O (nx5631z1), .CI (
          nx5630z1), .DI (conv_core_inst_for_i_sva[12]), .S (nx5630z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_17 (.O (nx5632z1), .CI (
          nx5631z1), .DI (conv_core_inst_for_i_sva[13]), .S (nx5631z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_18 (.O (nx5633z1), .CI (
          nx5632z1), .DI (conv_core_inst_for_i_sva[14]), .S (nx5632z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_19 (.O (nx6621z1), .CI (
          nx5633z1), .DI (conv_core_inst_for_i_sva[15]), .S (nx5633z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_20 (.O (nx6622z1), .CI (
          nx6621z1), .DI (conv_core_inst_for_i_sva[16]), .S (nx6621z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_21 (.O (nx6623z1), .CI (
          nx6622z1), .DI (conv_core_inst_for_i_sva[17]), .S (nx6622z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_22 (.O (nx6624z1), .CI (
          nx6623z1), .DI (conv_core_inst_for_i_sva[18]), .S (nx6623z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_23 (.O (nx6625z1), .CI (
          nx6624z1), .DI (conv_core_inst_for_i_sva[19]), .S (nx6624z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_24 (.O (nx6626z1), .CI (
          nx6625z1), .DI (conv_core_inst_for_i_sva[20]), .S (nx6625z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_25 (.O (nx6627z1), .CI (
          nx6626z1), .DI (conv_core_inst_for_i_sva[21]), .S (nx6626z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_26 (.O (nx6628z1), .CI (
          nx6627z1), .DI (conv_core_inst_for_i_sva[22]), .S (nx6627z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_27 (.O (nx6629z1), .CI (
          nx6628z1), .DI (conv_core_inst_for_i_sva[23]), .S (nx6628z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_28 (.O (nx6630z1), .CI (
          nx6629z1), .DI (conv_core_inst_for_i_sva[24]), .S (nx6629z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_29 (.O (nx7618z1), .CI (
          nx6630z1), .DI (conv_core_inst_for_i_sva[25]), .S (nx6630z2)) ;
    MUXCY for_for_for_for_acc_3_tmp_add32_3_muxcy_30 (.O (nx7619z1), .CI (
          nx7618z1), .DI (conv_core_inst_for_i_sva[26]), .S (nx7618z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_0 (.O (nx34916z1), .CI (px1140), .DI (
          \z_out_4(0)  ), .S (nx34917z1)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_1 (.O (nx34915z1), .CI (nx34916z1), .DI (
          \z_out_4(1)  ), .S (nx34916z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_2 (.O (nx34914z1), .CI (nx34915z1), .DI (
          \z_out_4(2)  ), .S (nx34915z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_3 (.O (nx34913z1), .CI (nx34914z1), .DI (
          \z_out_4(3)  ), .S (nx34914z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_4 (.O (nx34912z1), .CI (nx34913z1), .DI (
          \z_out_4(4)  ), .S (nx34913z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_5 (.O (nx34911z1), .CI (nx34912z1), .DI (
          \z_out_4(5)  ), .S (nx34912z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_6 (.O (nx34910z1), .CI (nx34911z1), .DI (
          \z_out_4(6)  ), .S (nx34911z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_7 (.O (nx34909z1), .CI (nx34910z1), .DI (
          \z_out_4(7)  ), .S (nx34910z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_8 (.O (nx34908z1), .CI (nx34909z1), .DI (
          \z_out_4(8)  ), .S (nx34909z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_9 (.O (nx53948z1), .CI (nx34908z1), .DI (
          \z_out_4(9)  ), .S (nx34908z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_10 (.O (nx53949z1), .CI (nx53948z1), .DI (
          \z_out_4(10)  ), .S (nx53948z2)) ;
    MUXCY image_rsci_addr_d_add13_4_muxcy_11 (.O (nx38873z1), .CI (nx53949z1), .DI (
          \z_out_4(11)  ), .S (nx53949z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_0 (.O (nx34262z1), .CI (
          px1551), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[0]), .S (
          nx34261z1)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_1 (.O (nx34263z1), .CI (
          nx34262z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[1]), .S (
          nx34262z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_2 (.O (nx34264z1), .CI (
          nx34263z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[2]), .S (
          nx34263z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_3 (.O (nx34265z1), .CI (
          nx34264z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[3]), .S (
          nx34264z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_4 (.O (nx34266z1), .CI (
          nx34265z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[4]), .S (
          nx34265z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_5 (.O (nx34267z1), .CI (
          nx34266z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[5]), .S (
          nx34266z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_6 (.O (nx34268z1), .CI (
          nx34267z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[6]), .S (
          nx34267z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_7 (.O (nx34269z1), .CI (
          nx34268z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[7]), .S (
          nx34268z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_8 (.O (nx34270z1), .CI (
          nx34269z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[8]), .S (
          nx34269z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_9 (.O (nx50530z1), .CI (
          nx34270z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[9]), .S (
          nx34270z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_10 (.O (nx50529z1), .CI (
          nx50530z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[10]), .S (
          nx50530z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_11 (.O (nx50528z1), .CI (
          nx50529z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[11]), .S (
          nx50529z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_12 (.O (nx50527z1), .CI (
          nx50528z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[12]), .S (
          nx50528z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_13 (.O (nx50526z1), .CI (
          nx50527z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[13]), .S (
          nx50527z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_14 (.O (nx50525z1), .CI (
          nx50526z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[14]), .S (
          nx50526z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_15 (.O (nx50524z1), .CI (
          nx50525z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[15]), .S (
          nx50525z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_16 (.O (nx50523z1), .CI (
          nx50524z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[16]), .S (
          nx50524z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_17 (.O (nx50522z1), .CI (
          nx50523z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[17]), .S (
          nx50523z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_18 (.O (nx50521z1), .CI (
          nx50522z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[18]), .S (
          nx50522z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_19 (.O (nx49533z1), .CI (
          nx50521z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[19]), .S (
          nx50521z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_20 (.O (nx49532z1), .CI (
          nx49533z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[20]), .S (
          nx49533z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_21 (.O (nx49531z1), .CI (
          nx49532z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[21]), .S (
          nx49532z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_22 (.O (nx49530z1), .CI (
          nx49531z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[22]), .S (
          nx49531z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_23 (.O (nx49529z1), .CI (
          nx49530z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[23]), .S (
          nx49530z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_24 (.O (nx49528z1), .CI (
          nx49529z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[24]), .S (
          nx49529z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_25 (.O (nx49527z1), .CI (
          nx49528z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[25]), .S (
          nx49528z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_26 (.O (nx49526z1), .CI (
          nx49527z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[26]), .S (
          nx49527z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_27 (.O (nx49525z1), .CI (
          nx49526z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[27]), .S (
          nx49526z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_28 (.O (nx49524z1), .CI (
          nx49525z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[28]), .S (
          nx49525z2)) ;
    MUXCY for_for_for_for_aif_acc_nl_sub31_11_muxcy_29 (.O (nx48536z1), .CI (
          nx49524z1), .DI (conv_core_inst_for_for_for_for_acc_3_tmp[29]), .S (
          nx49524z2)) ;
    MUXCY muxcy_0_1 (.O (nx39518z1), .CI (nx39517z1), .DI (nx39517z2), .S (
          nx39517z5)) ;
    MUXCY muxcy_0_2 (.O (nx39519z1), .CI (nx39518z1), .DI (nx39518z2), .S (
          nx39518z3)) ;
    MUXCY muxcy_0_3 (.O (nx39520z1), .CI (nx39519z1), .DI (nx39519z2), .S (
          nx39519z3)) ;
    MUXCY muxcy_0_4 (.O (nx39521z1), .CI (nx39520z1), .DI (nx39520z2), .S (
          nx39520z3)) ;
    MUXCY muxcy_0_5 (.O (nx39522z1), .CI (nx39521z1), .DI (nx39521z2), .S (
          nx39521z3)) ;
    MUXCY muxcy_0_6 (.O (nx39523z1), .CI (nx39522z1), .DI (nx39522z2), .S (
          nx39522z3)) ;
    MUXCY muxcy_0_7 (.O (nx50037z1), .CI (nx39523z1), .DI (nx39523z2), .S (
          nx39523z3)) ;
    MUXCY z_out_1_add34_7_muxcy_0 (.O (nx28349z1), .CI (not_fsm_output_5), .DI (
          nx28350z1), .S (nx28350z3)) ;
    MUXCY z_out_1_add34_7_muxcy_1 (.O (nx28348z1), .CI (nx28349z1), .DI (
          nx28349z2), .S (nx28349z3)) ;
    MUXCY z_out_1_add34_7_muxcy_2 (.O (nx28347z1), .CI (nx28348z1), .DI (
          nx28348z2), .S (nx28348z3)) ;
    MUXCY z_out_1_add34_7_muxcy_3 (.O (nx28346z1), .CI (nx28347z1), .DI (
          nx28347z2), .S (nx28347z3)) ;
    MUXCY z_out_1_add34_7_muxcy_4 (.O (nx28345z1), .CI (nx28346z1), .DI (
          nx28346z2), .S (nx28346z3)) ;
    MUXCY z_out_1_add34_7_muxcy_5 (.O (nx28344z1), .CI (nx28345z1), .DI (
          nx28345z2), .S (nx28345z3)) ;
    MUXCY z_out_1_add34_7_muxcy_6 (.O (nx28343z1), .CI (nx28344z1), .DI (
          nx28344z2), .S (nx28344z3)) ;
    MUXCY z_out_1_add34_7_muxcy_7 (.O (nx28342z1), .CI (nx28343z1), .DI (
          nx28343z2), .S (nx28343z3)) ;
    MUXCY z_out_1_add34_7_muxcy_8 (.O (nx28341z1), .CI (nx28342z1), .DI (
          nx28342z2), .S (nx28342z3)) ;
    MUXCY z_out_1_add34_7_muxcy_9 (.O (nx47647z1), .CI (nx28341z1), .DI (
          nx28341z2), .S (nx28341z3)) ;
    MUXCY z_out_1_add34_7_muxcy_10 (.O (nx47648z1), .CI (nx47647z1), .DI (
          nx47647z2), .S (nx47647z3)) ;
    MUXCY z_out_1_add34_7_muxcy_11 (.O (nx47649z1), .CI (nx47648z1), .DI (
          nx47648z2), .S (nx47648z3)) ;
    MUXCY z_out_1_add34_7_muxcy_12 (.O (nx47650z1), .CI (nx47649z1), .DI (
          nx47649z2), .S (nx47649z3)) ;
    MUXCY z_out_1_add34_7_muxcy_13 (.O (nx47651z1), .CI (nx47650z1), .DI (
          nx47650z2), .S (nx47650z3)) ;
    MUXCY z_out_1_add34_7_muxcy_14 (.O (nx47652z1), .CI (nx47651z1), .DI (
          nx47651z2), .S (nx47651z3)) ;
    MUXCY z_out_1_add34_7_muxcy_15 (.O (nx47653z1), .CI (nx47652z1), .DI (
          nx47652z2), .S (nx47652z3)) ;
    MUXCY z_out_1_add34_7_muxcy_16 (.O (nx47654z2), .CI (nx47653z1), .DI (
          nx47653z2), .S (nx47653z3)) ;
    MUXCY z_out_1_add34_7_muxcy_17 (.O (nx47655z1), .CI (nx47654z2), .DI (
          nx47654z3), .S (nx47654z4)) ;
    MUXCY z_out_1_add34_7_muxcy_18 (.O (nx47656z1), .CI (nx47655z1), .DI (
          nx47655z2), .S (nx47655z3)) ;
    MUXCY z_out_1_add34_7_muxcy_19 (.O (nx48644z1), .CI (nx47656z1), .DI (
          nx47656z2), .S (nx47656z3)) ;
    MUXCY z_out_1_add34_7_muxcy_20 (.O (nx48645z1), .CI (nx48644z1), .DI (
          nx48644z2), .S (nx48644z3)) ;
    MUXCY z_out_1_add34_7_muxcy_21 (.O (nx48646z1), .CI (nx48645z1), .DI (
          nx48645z2), .S (nx48645z3)) ;
    MUXCY z_out_1_add34_7_muxcy_22 (.O (nx48647z1), .CI (nx48646z1), .DI (
          nx48646z2), .S (nx48646z3)) ;
    MUXCY z_out_1_add34_7_muxcy_23 (.O (nx48648z1), .CI (nx48647z1), .DI (
          nx48647z2), .S (nx48647z3)) ;
    MUXCY z_out_1_add34_7_muxcy_24 (.O (nx48649z1), .CI (nx48648z1), .DI (
          nx48648z2), .S (nx48648z3)) ;
    MUXCY z_out_1_add34_7_muxcy_25 (.O (nx48650z1), .CI (nx48649z1), .DI (
          nx48649z2), .S (nx48649z3)) ;
    MUXCY z_out_1_add34_7_muxcy_26 (.O (nx48651z2), .CI (nx48650z1), .DI (
          nx48650z2), .S (nx48650z3)) ;
    MUXCY z_out_1_add34_7_muxcy_27 (.O (nx48652z1), .CI (nx48651z2), .DI (
          nx48651z3), .S (nx48651z4)) ;
    MUXCY z_out_1_add34_7_muxcy_28 (.O (nx48653z1), .CI (nx48652z1), .DI (
          nx48652z2), .S (nx48652z3)) ;
    MUXCY z_out_1_add34_7_muxcy_29 (.O (nx49641z1), .CI (nx48653z1), .DI (
          nx48653z2), .S (nx48653z3)) ;
    MUXCY z_out_1_add34_7_muxcy_30 (.O (nx49642z1), .CI (nx49641z1), .DI (
          nx49641z2), .S (nx49641z3)) ;
    MUXCY z_out_1_add34_7_muxcy_31 (.O (nx34566z1), .CI (nx49642z1), .DI (
          nx49642z2), .S (nx49642z4)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(31)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[0]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[0]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(30)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[1]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[1]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(29)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[2]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[2]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(28)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[3]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[3]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(27)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[4]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[4]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(26)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[5]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[5]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(25)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[6]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[6]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(24)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[7]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[7]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(23)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[8]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[8]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(22)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[9]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[9]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(21)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[10]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[10]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(20)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[11]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[11]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(19)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[12]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[12]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(18)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[13]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[13]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(17)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[14]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[14]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(16)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[15]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[15]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(15)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[16]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[16]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(14)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[17]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[17]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(13)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[18]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[18]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(12)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[19]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[19]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(11)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[20]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[20]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(10)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[21]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[21]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(9)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[22]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[22]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(8)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[23]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[23]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(7)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[24]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[24]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(6)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[25]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[25]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(5)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[26]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[26]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(4)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[27]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[27]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(3)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[28]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[28]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(2)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[29]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[29]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(1)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[30]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[30]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_7_itm_2(0)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_7_itm_2[31]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_sortie_rsc_data_out_int[31]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(31)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[0]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[0]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(30)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[1]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[1]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(29)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[2]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[2]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(28)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[3]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[3]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(27)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[4]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[4]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(26)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[5]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[5]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(25)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[6]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[6]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(24)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[7]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[7]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(23)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[8]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[8]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(22)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[9]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[9]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(21)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[10]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[10]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(20)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[11]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[11]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(19)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[12]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[12]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(18)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[13]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[13]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(17)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[14]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[14]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(16)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[15]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[15]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(15)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[16]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[16]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(14)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[17]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[17]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(13)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[18]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[18]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(12)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[19]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[19]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(11)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[20]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[20]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(10)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[21]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[21]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(9)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[22]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[22]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(8)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[23]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[23]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(7)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[24]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[24]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(6)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[25]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[25]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(5)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[26]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[26]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(4)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[27]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[27]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(3)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[28]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[28]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(2)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[29]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[29]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(1)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[30]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[30]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_asn_6_itm_2(0)  (.Q (
         conv_core_inst_for_for_for_for_if_asn_6_itm_2[31]), .C (p_clk_int), .CE (
         nx39517z3), .D (p_nbus_kernel_rsc_data_out_int[31]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(12)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[0]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[12]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(11)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[1]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[11]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(10)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[2]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[10]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(9)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[3]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[9]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(8)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[4]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[8]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(7)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[5]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[7]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(6)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[6]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[6]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(5)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[7]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[5]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(4)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[8]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[4]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(3)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[9]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[3]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(2)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[10]), .C (p_clk_int
         ), .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[2]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(1)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[11]), .C (p_clk_int
         ), .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[1]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_ii_28_0_itm_2(0)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_ii_28_0_itm_2[12]), .C (p_clk_int
         ), .CE (nx39517z3), .D (conv_core_inst_for_for_for_for_acc_3_tmp[0]), .R (
         p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(12)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[0]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[15]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(11)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[1]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[14]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(10)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[2]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[13]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(9)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[3]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[12]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(8)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[4]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[11]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(7)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[5]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[10]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(6)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[6]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[9]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(5)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[7]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[8]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(4)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[8]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[7]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(3)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[9]), .C (p_clk_int)
         , .CE (nx39517z3), .D (conv_core_inst_jj_sva[6]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(2)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[10]), .C (p_clk_int
         ), .CE (nx39517z3), .D (conv_core_inst_jj_sva[5]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(1)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[11]), .C (p_clk_int
         ), .CE (nx39517z3), .D (conv_core_inst_jj_sva[4]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_15_3_itm_2(0)  (.Q (
         conv_core_inst_for_for_for_for_if_slc_jj_15_3_itm_2[12]), .C (p_clk_int
         ), .CE (nx39517z3), .D (conv_core_inst_jj_sva[3]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_2_0_itm_3(2)  (.Q (
         p_nbus_image_rsc_addr_1_0[13]), .C (p_clk_int), .CE (nx39517z3), .D (
         conv_core_inst_jj_sva[2]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_2_0_itm_3(1)  (.Q (
         p_nbus_image_rsc_addr_1_0[14]), .C (p_clk_int), .CE (nx39517z3), .D (
         conv_core_inst_jj_sva[1]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_if_slc_jj_2_0_itm_3(0)  (.Q (
         p_nbus_image_rsc_addr_1_0[15]), .C (p_clk_int), .CE (nx39517z3), .D (
         conv_core_inst_jj_sva[0]), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva(4)  (.Q (\for_for_for_for_n_4_0_sva(4)  
         ), .C (p_clk_int), .CE (nx39517z3), .D (nx1713z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva(3)  (.Q (
         conv_core_inst_for_for_for_for_n_4_0_sva[4]), .C (p_clk_int), .CE (
         nx39517z3), .D (nx2710z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva(2)  (.Q (\for_for_for_for_n_4_0_sva(2)  
         ), .C (p_clk_int), .CE (nx39517z3), .D (nx3707z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva(1)  (.Q (\for_for_for_for_n_4_0_sva(1)  
         ), .C (p_clk_int), .CE (nx39517z3), .D (nx4704z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_for_for_n_4_0_sva(0)  (.Q (\for_for_for_for_n_4_0_sva(0)  
         ), .C (p_clk_int), .CE (nx39517z3), .D (nx5701z1), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(9)  (.Q (\p_fsm_output(10)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (nx22387z1), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(8)  (.Q (\fsm_output(9)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (nx21390z1), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(7)  (.Q (\fsm_output(8)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (nx20393z1), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(6)  (.Q (\fsm_output(7)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (nx19396z1), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(5)  (.Q (\fsm_output(6)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (\fsm_output(5)  ), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(4)  (.Q (\fsm_output(5)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (\fsm_output(4)  ), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(3)  (.Q (\fsm_output(4)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (\fsm_output(3)  ), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(2)  (.Q (\fsm_output(3)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (nx15408z1), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(1)  (.Q (
         \conv_core_core_fsm_inst_fsm_output(2)  ), .C (p_clk_int), .CE (
         nx39517z3), .D (nx14411z1), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(0)  (.Q (\fsm_output(1)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (nx13414z1), .R (p_rst_int)) ;
    FDRE \conv_core_core_fsm_inst_reg_state_var(10)  (.Q (\fsm_output(0)  ), .C (
         p_clk_int), .CE (nx39517z3), .D (nx43133z1), .R (nx39517z1)) ;
endmodule


module inc_31_0 ( cin, a, d, cout, \p_rows_rsc_z_int(30)  , \p_fsm_output(9)  , 
                  \p_fsm_output(0)  , \p_for_i_sva(30)  , px1533, 
                  \p_rows_rsc_z_int(29)  , \p_for_i_sva(29)  , px1531, 
                  \p_rows_rsc_z_int(28)  , \p_for_i_sva(28)  , px1529, 
                  \p_rows_rsc_z_int(27)  , \p_for_i_sva(27)  , px1527, 
                  \p_rows_rsc_z_int(26)  , \p_for_i_sva(26)  , px1525, 
                  \p_rows_rsc_z_int(25)  , \p_for_i_sva(25)  , px1523, 
                  \p_rows_rsc_z_int(24)  , \p_for_i_sva(24)  , px1521, 
                  \p_rows_rsc_z_int(23)  , \p_for_i_sva(23)  , px1519, 
                  \p_rows_rsc_z_int(22)  , \p_for_i_sva(22)  , px1517, 
                  \p_rows_rsc_z_int(21)  , \p_for_i_sva(21)  , px1515, 
                  \p_rows_rsc_z_int(20)  , \p_for_i_sva(20)  , px1513, 
                  \p_rows_rsc_z_int(19)  , \p_for_i_sva(19)  , px1511, 
                  \p_rows_rsc_z_int(18)  , \p_for_i_sva(18)  , px1509, 
                  \p_rows_rsc_z_int(17)  , \p_for_i_sva(17)  , px1507, 
                  \p_rows_rsc_z_int(16)  , \p_for_i_sva(16)  , px1505, 
                  \p_rows_rsc_z_int(15)  , \p_for_i_sva(15)  , px1503, 
                  \p_rows_rsc_z_int(14)  , \p_for_i_sva(14)  , px1501, 
                  \p_rows_rsc_z_int(13)  , \p_for_i_sva(13)  , px1499, 
                  \p_rows_rsc_z_int(12)  , \p_for_i_sva(12)  , px1497, 
                  \p_rows_rsc_z_int(11)  , \p_for_i_sva(11)  , px1495, 
                  \p_rows_rsc_z_int(10)  , \p_for_i_sva(10)  , px1493, 
                  \p_rows_rsc_z_int(9)  , \p_for_i_sva(9)  , px1491, 
                  \p_rows_rsc_z_int(8)  , \p_for_i_sva(8)  , px1489, 
                  \p_rows_rsc_z_int(7)  , \p_for_i_sva(7)  , px1487, 
                  \p_rows_rsc_z_int(6)  , \p_for_i_sva(6)  , px1485, 
                  \p_rows_rsc_z_int(5)  , \p_for_i_sva(5)  , px1483, 
                  \p_rows_rsc_z_int(4)  , \p_for_i_sva(4)  , px1481, 
                  \p_rows_rsc_z_int(3)  , \p_for_i_sva(3)  , px1479, 
                  \p_sortie_rsc_addr_1_0(2)  , \p_rows_rsc_z_int(2)  , 
                  \p_fsm_output(8)  , px1477, \p_sortie_rsc_addr_1_0(1)  , 
                  \p_rows_rsc_z_int(1)  , px1475, \p_sortie_rsc_addr_1_0(0)  , 
                  \p_rows_rsc_z_int(0)  , px1473 ) ;

    input cin ;
    input [30:0]a ;
    output [30:0]d ;
    output cout ;
    input \p_rows_rsc_z_int(30)   ;
    input \p_fsm_output(9)   ;
    input \p_fsm_output(0)   ;
    input \p_for_i_sva(30)   ;
    input px1533 ;
    input \p_rows_rsc_z_int(29)   ;
    input \p_for_i_sva(29)   ;
    input px1531 ;
    input \p_rows_rsc_z_int(28)   ;
    input \p_for_i_sva(28)   ;
    input px1529 ;
    input \p_rows_rsc_z_int(27)   ;
    input \p_for_i_sva(27)   ;
    input px1527 ;
    input \p_rows_rsc_z_int(26)   ;
    input \p_for_i_sva(26)   ;
    input px1525 ;
    input \p_rows_rsc_z_int(25)   ;
    input \p_for_i_sva(25)   ;
    input px1523 ;
    input \p_rows_rsc_z_int(24)   ;
    input \p_for_i_sva(24)   ;
    input px1521 ;
    input \p_rows_rsc_z_int(23)   ;
    input \p_for_i_sva(23)   ;
    input px1519 ;
    input \p_rows_rsc_z_int(22)   ;
    input \p_for_i_sva(22)   ;
    input px1517 ;
    input \p_rows_rsc_z_int(21)   ;
    input \p_for_i_sva(21)   ;
    input px1515 ;
    input \p_rows_rsc_z_int(20)   ;
    input \p_for_i_sva(20)   ;
    input px1513 ;
    input \p_rows_rsc_z_int(19)   ;
    input \p_for_i_sva(19)   ;
    input px1511 ;
    input \p_rows_rsc_z_int(18)   ;
    input \p_for_i_sva(18)   ;
    input px1509 ;
    input \p_rows_rsc_z_int(17)   ;
    input \p_for_i_sva(17)   ;
    input px1507 ;
    input \p_rows_rsc_z_int(16)   ;
    input \p_for_i_sva(16)   ;
    input px1505 ;
    input \p_rows_rsc_z_int(15)   ;
    input \p_for_i_sva(15)   ;
    input px1503 ;
    input \p_rows_rsc_z_int(14)   ;
    input \p_for_i_sva(14)   ;
    input px1501 ;
    input \p_rows_rsc_z_int(13)   ;
    input \p_for_i_sva(13)   ;
    input px1499 ;
    input \p_rows_rsc_z_int(12)   ;
    input \p_for_i_sva(12)   ;
    input px1497 ;
    input \p_rows_rsc_z_int(11)   ;
    input \p_for_i_sva(11)   ;
    input px1495 ;
    input \p_rows_rsc_z_int(10)   ;
    input \p_for_i_sva(10)   ;
    input px1493 ;
    input \p_rows_rsc_z_int(9)   ;
    input \p_for_i_sva(9)   ;
    input px1491 ;
    input \p_rows_rsc_z_int(8)   ;
    input \p_for_i_sva(8)   ;
    input px1489 ;
    input \p_rows_rsc_z_int(7)   ;
    input \p_for_i_sva(7)   ;
    input px1487 ;
    input \p_rows_rsc_z_int(6)   ;
    input \p_for_i_sva(6)   ;
    input px1485 ;
    input \p_rows_rsc_z_int(5)   ;
    input \p_for_i_sva(5)   ;
    input px1483 ;
    input \p_rows_rsc_z_int(4)   ;
    input \p_for_i_sva(4)   ;
    input px1481 ;
    input \p_rows_rsc_z_int(3)   ;
    input \p_for_i_sva(3)   ;
    input px1479 ;
    input \p_sortie_rsc_addr_1_0(2)   ;
    input \p_rows_rsc_z_int(2)   ;
    input \p_fsm_output(8)   ;
    input px1477 ;
    input \p_sortie_rsc_addr_1_0(1)   ;
    input \p_rows_rsc_z_int(1)   ;
    input px1475 ;
    input \p_sortie_rsc_addr_1_0(0)   ;
    input \p_rows_rsc_z_int(0)   ;
    input px1473 ;

    wire nx8473z2, nx8473z1, nx8473z3, nx8474z1, nx8474z2, nx8475z1, nx8475z2, 
         nx8476z1, nx8476z2, nx8477z1, nx8477z2, nx8478z1, nx8478z2, nx8479z1, 
         nx8479z2, nx8480z1, nx8480z2, nx8481z1, nx8481z2, nx8482z1, nx8482z2, 
         nx60018z1, nx60018z2, nx60019z1, nx60019z2, nx60020z1, nx60020z2, 
         nx60021z1, nx60021z2, nx60022z1, nx60022z2, nx60023z1, nx60023z2, 
         nx60024z1, nx60024z2, nx60025z1, nx60025z2, nx60026z1, nx60026z2, 
         nx60027z1, nx60027z2, nx61015z1, nx61015z2, nx61016z1, nx61016z2, 
         nx61017z1, nx61017z2, nx61018z1, nx61018z2, nx61019z1, nx61019z2, 
         nx61020z1, nx61020z2, nx61021z1, nx61021z2, nx61022z1, nx61022z2, 
         nx61023z1, nx61023z2, nx61024z1, nx61024z2, nx18601z1, nx18601z2;



    GND ps_gnd (.G (nx8473z2)) ;
    VCC ps_vcc (.P (nx8473z1)) ;
    XORCY xorcy_0 (.O (d[0]), .CI (nx8473z1), .LI (nx8473z3)) ;
    XORCY xorcy_1 (.O (d[1]), .CI (nx8474z1), .LI (nx8474z2)) ;
    XORCY xorcy_2 (.O (d[2]), .CI (nx8475z1), .LI (nx8475z2)) ;
    XORCY xorcy_3 (.O (d[3]), .CI (nx8476z1), .LI (nx8476z2)) ;
    XORCY xorcy_4 (.O (d[4]), .CI (nx8477z1), .LI (nx8477z2)) ;
    XORCY xorcy_5 (.O (d[5]), .CI (nx8478z1), .LI (nx8478z2)) ;
    XORCY xorcy_6 (.O (d[6]), .CI (nx8479z1), .LI (nx8479z2)) ;
    XORCY xorcy_7 (.O (d[7]), .CI (nx8480z1), .LI (nx8480z2)) ;
    XORCY xorcy_8 (.O (d[8]), .CI (nx8481z1), .LI (nx8481z2)) ;
    XORCY xorcy_9 (.O (d[9]), .CI (nx8482z1), .LI (nx8482z2)) ;
    XORCY xorcy_10 (.O (d[10]), .CI (nx60018z1), .LI (nx60018z2)) ;
    XORCY xorcy_11 (.O (d[11]), .CI (nx60019z1), .LI (nx60019z2)) ;
    XORCY xorcy_12 (.O (d[12]), .CI (nx60020z1), .LI (nx60020z2)) ;
    XORCY xorcy_13 (.O (d[13]), .CI (nx60021z1), .LI (nx60021z2)) ;
    XORCY xorcy_14 (.O (d[14]), .CI (nx60022z1), .LI (nx60022z2)) ;
    XORCY xorcy_15 (.O (d[15]), .CI (nx60023z1), .LI (nx60023z2)) ;
    XORCY xorcy_16 (.O (d[16]), .CI (nx60024z1), .LI (nx60024z2)) ;
    XORCY xorcy_17 (.O (d[17]), .CI (nx60025z1), .LI (nx60025z2)) ;
    XORCY xorcy_18 (.O (d[18]), .CI (nx60026z1), .LI (nx60026z2)) ;
    XORCY xorcy_19 (.O (d[19]), .CI (nx60027z1), .LI (nx60027z2)) ;
    XORCY xorcy_20 (.O (d[20]), .CI (nx61015z1), .LI (nx61015z2)) ;
    XORCY xorcy_21 (.O (d[21]), .CI (nx61016z1), .LI (nx61016z2)) ;
    XORCY xorcy_22 (.O (d[22]), .CI (nx61017z1), .LI (nx61017z2)) ;
    XORCY xorcy_23 (.O (d[23]), .CI (nx61018z1), .LI (nx61018z2)) ;
    XORCY xorcy_24 (.O (d[24]), .CI (nx61019z1), .LI (nx61019z2)) ;
    XORCY xorcy_25 (.O (d[25]), .CI (nx61020z1), .LI (nx61020z2)) ;
    XORCY xorcy_26 (.O (d[26]), .CI (nx61021z1), .LI (nx61021z2)) ;
    XORCY xorcy_27 (.O (d[27]), .CI (nx61022z1), .LI (nx61022z2)) ;
    XORCY xorcy_28 (.O (d[28]), .CI (nx61023z1), .LI (nx61023z2)) ;
    XORCY xorcy_29 (.O (d[29]), .CI (nx61024z1), .LI (nx61024z2)) ;
    XORCY xorcy_30 (.O (d[30]), .CI (nx18601z1), .LI (nx18601z2)) ;
    MUXCY muxcy_30 (.O (cout), .CI (nx18601z1), .DI (nx8473z2), .S (nx18601z2)
          ) ;
    MUXCY muxcy_0 (.O (nx8474z1), .CI (nx8473z1), .DI (nx8473z2), .S (nx8473z3)
          ) ;
    MUXCY muxcy_1 (.O (nx8475z1), .CI (nx8474z1), .DI (nx8473z2), .S (nx8474z2)
          ) ;
    MUXCY muxcy_2 (.O (nx8476z1), .CI (nx8475z1), .DI (nx8473z2), .S (nx8475z2)
          ) ;
    MUXCY muxcy_3 (.O (nx8477z1), .CI (nx8476z1), .DI (nx8473z2), .S (nx8476z2)
          ) ;
    MUXCY muxcy_4 (.O (nx8478z1), .CI (nx8477z1), .DI (nx8473z2), .S (nx8477z2)
          ) ;
    MUXCY muxcy_5 (.O (nx8479z1), .CI (nx8478z1), .DI (nx8473z2), .S (nx8478z2)
          ) ;
    MUXCY muxcy_6 (.O (nx8480z1), .CI (nx8479z1), .DI (nx8473z2), .S (nx8479z2)
          ) ;
    MUXCY muxcy_7 (.O (nx8481z1), .CI (nx8480z1), .DI (nx8473z2), .S (nx8480z2)
          ) ;
    MUXCY muxcy_8 (.O (nx8482z1), .CI (nx8481z1), .DI (nx8473z2), .S (nx8481z2)
          ) ;
    MUXCY muxcy_9 (.O (nx60018z1), .CI (nx8482z1), .DI (nx8473z2), .S (nx8482z2)
          ) ;
    MUXCY muxcy_10 (.O (nx60019z1), .CI (nx60018z1), .DI (nx8473z2), .S (
          nx60018z2)) ;
    MUXCY muxcy_11 (.O (nx60020z1), .CI (nx60019z1), .DI (nx8473z2), .S (
          nx60019z2)) ;
    MUXCY muxcy_12 (.O (nx60021z1), .CI (nx60020z1), .DI (nx8473z2), .S (
          nx60020z2)) ;
    MUXCY muxcy_13 (.O (nx60022z1), .CI (nx60021z1), .DI (nx8473z2), .S (
          nx60021z2)) ;
    MUXCY muxcy_14 (.O (nx60023z1), .CI (nx60022z1), .DI (nx8473z2), .S (
          nx60022z2)) ;
    MUXCY muxcy_15 (.O (nx60024z1), .CI (nx60023z1), .DI (nx8473z2), .S (
          nx60023z2)) ;
    MUXCY muxcy_16 (.O (nx60025z1), .CI (nx60024z1), .DI (nx8473z2), .S (
          nx60024z2)) ;
    MUXCY muxcy_17 (.O (nx60026z1), .CI (nx60025z1), .DI (nx8473z2), .S (
          nx60025z2)) ;
    MUXCY muxcy_18 (.O (nx60027z1), .CI (nx60026z1), .DI (nx8473z2), .S (
          nx60026z2)) ;
    MUXCY muxcy_19 (.O (nx61015z1), .CI (nx60027z1), .DI (nx8473z2), .S (
          nx60027z2)) ;
    MUXCY muxcy_20 (.O (nx61016z1), .CI (nx61015z1), .DI (nx8473z2), .S (
          nx61015z2)) ;
    MUXCY muxcy_21 (.O (nx61017z1), .CI (nx61016z1), .DI (nx8473z2), .S (
          nx61016z2)) ;
    MUXCY muxcy_22 (.O (nx61018z1), .CI (nx61017z1), .DI (nx8473z2), .S (
          nx61017z2)) ;
    MUXCY muxcy_23 (.O (nx61019z1), .CI (nx61018z1), .DI (nx8473z2), .S (
          nx61018z2)) ;
    MUXCY muxcy_24 (.O (nx61020z1), .CI (nx61019z1), .DI (nx8473z2), .S (
          nx61019z2)) ;
    MUXCY muxcy_25 (.O (nx61021z1), .CI (nx61020z1), .DI (nx8473z2), .S (
          nx61020z2)) ;
    MUXCY muxcy_26 (.O (nx61022z1), .CI (nx61021z1), .DI (nx8473z2), .S (
          nx61021z2)) ;
    MUXCY muxcy_27 (.O (nx61023z1), .CI (nx61022z1), .DI (nx8473z2), .S (
          nx61022z2)) ;
    MUXCY muxcy_28 (.O (nx61024z1), .CI (nx61023z1), .DI (nx8473z2), .S (
          nx61023z2)) ;
    MUXCY muxcy_29 (.O (nx18601z1), .CI (nx61024z1), .DI (nx8473z2), .S (
          nx61024z2)) ;
    LUT5 ix18601z1313 (.O (nx18601z2), .I0 (\p_rows_rsc_z_int(30)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(30)  )
         , .I4 (px1533)) ;
         defparam ix18601z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61024z1313 (.O (nx61024z2), .I0 (\p_rows_rsc_z_int(29)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(29)  )
         , .I4 (px1531)) ;
         defparam ix61024z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61023z1313 (.O (nx61023z2), .I0 (\p_rows_rsc_z_int(28)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(28)  )
         , .I4 (px1529)) ;
         defparam ix61023z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61022z1313 (.O (nx61022z2), .I0 (\p_rows_rsc_z_int(27)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(27)  )
         , .I4 (px1527)) ;
         defparam ix61022z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61021z1313 (.O (nx61021z2), .I0 (\p_rows_rsc_z_int(26)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(26)  )
         , .I4 (px1525)) ;
         defparam ix61021z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61020z1313 (.O (nx61020z2), .I0 (\p_rows_rsc_z_int(25)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(25)  )
         , .I4 (px1523)) ;
         defparam ix61020z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61019z1313 (.O (nx61019z2), .I0 (\p_rows_rsc_z_int(24)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(24)  )
         , .I4 (px1521)) ;
         defparam ix61019z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61018z1313 (.O (nx61018z2), .I0 (\p_rows_rsc_z_int(23)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(23)  )
         , .I4 (px1519)) ;
         defparam ix61018z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61017z1313 (.O (nx61017z2), .I0 (\p_rows_rsc_z_int(22)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(22)  )
         , .I4 (px1517)) ;
         defparam ix61017z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61016z1313 (.O (nx61016z2), .I0 (\p_rows_rsc_z_int(21)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(21)  )
         , .I4 (px1515)) ;
         defparam ix61016z1313.INIT = 32'hDC50FFFF;
    LUT5 ix61015z1313 (.O (nx61015z2), .I0 (\p_rows_rsc_z_int(20)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(20)  )
         , .I4 (px1513)) ;
         defparam ix61015z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60027z1313 (.O (nx60027z2), .I0 (\p_rows_rsc_z_int(19)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(19)  )
         , .I4 (px1511)) ;
         defparam ix60027z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60026z1313 (.O (nx60026z2), .I0 (\p_rows_rsc_z_int(18)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(18)  )
         , .I4 (px1509)) ;
         defparam ix60026z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60025z1313 (.O (nx60025z2), .I0 (\p_rows_rsc_z_int(17)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(17)  )
         , .I4 (px1507)) ;
         defparam ix60025z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60024z1313 (.O (nx60024z2), .I0 (\p_rows_rsc_z_int(16)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(16)  )
         , .I4 (px1505)) ;
         defparam ix60024z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60023z1313 (.O (nx60023z2), .I0 (\p_rows_rsc_z_int(15)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(15)  )
         , .I4 (px1503)) ;
         defparam ix60023z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60022z1313 (.O (nx60022z2), .I0 (\p_rows_rsc_z_int(14)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(14)  )
         , .I4 (px1501)) ;
         defparam ix60022z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60021z1313 (.O (nx60021z2), .I0 (\p_rows_rsc_z_int(13)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(13)  )
         , .I4 (px1499)) ;
         defparam ix60021z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60020z1313 (.O (nx60020z2), .I0 (\p_rows_rsc_z_int(12)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(12)  )
         , .I4 (px1497)) ;
         defparam ix60020z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60019z1313 (.O (nx60019z2), .I0 (\p_rows_rsc_z_int(11)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(11)  )
         , .I4 (px1495)) ;
         defparam ix60019z1313.INIT = 32'hDC50FFFF;
    LUT5 ix60018z1313 (.O (nx60018z2), .I0 (\p_rows_rsc_z_int(10)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(10)  )
         , .I4 (px1493)) ;
         defparam ix60018z1313.INIT = 32'hDC50FFFF;
    LUT5 ix8482z1313 (.O (nx8482z2), .I0 (\p_rows_rsc_z_int(9)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(9)  )
         , .I4 (px1491)) ;
         defparam ix8482z1313.INIT = 32'hDC50FFFF;
    LUT5 ix8481z1313 (.O (nx8481z2), .I0 (\p_rows_rsc_z_int(8)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(8)  )
         , .I4 (px1489)) ;
         defparam ix8481z1313.INIT = 32'hDC50FFFF;
    LUT5 ix8480z1313 (.O (nx8480z2), .I0 (\p_rows_rsc_z_int(7)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(7)  )
         , .I4 (px1487)) ;
         defparam ix8480z1313.INIT = 32'hDC50FFFF;
    LUT5 ix8479z1313 (.O (nx8479z2), .I0 (\p_rows_rsc_z_int(6)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(6)  )
         , .I4 (px1485)) ;
         defparam ix8479z1313.INIT = 32'hDC50FFFF;
    LUT5 ix8478z1313 (.O (nx8478z2), .I0 (\p_rows_rsc_z_int(5)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(5)  )
         , .I4 (px1483)) ;
         defparam ix8478z1313.INIT = 32'hDC50FFFF;
    LUT5 ix8477z1313 (.O (nx8477z2), .I0 (\p_rows_rsc_z_int(4)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(4)  )
         , .I4 (px1481)) ;
         defparam ix8477z1313.INIT = 32'hDC50FFFF;
    LUT5 ix8476z1313 (.O (nx8476z2), .I0 (\p_rows_rsc_z_int(3)  ), .I1 (
         \p_fsm_output(9)  ), .I2 (\p_fsm_output(0)  ), .I3 (\p_for_i_sva(3)  )
         , .I4 (px1479)) ;
         defparam ix8476z1313.INIT = 32'hDC50FFFF;
    LUT5 ix8475z1313 (.O (nx8475z2), .I0 (\p_sortie_rsc_addr_1_0(2)  ), .I1 (
         \p_rows_rsc_z_int(2)  ), .I2 (\p_fsm_output(8)  ), .I3 (
         \p_fsm_output(0)  ), .I4 (px1477)) ;
         defparam ix8475z1313.INIT = 32'hB3A0FFFF;
    LUT5 ix8474z1313 (.O (nx8474z2), .I0 (\p_sortie_rsc_addr_1_0(1)  ), .I1 (
         \p_rows_rsc_z_int(1)  ), .I2 (\p_fsm_output(8)  ), .I3 (
         \p_fsm_output(0)  ), .I4 (px1475)) ;
         defparam ix8474z1313.INIT = 32'hB3A0FFFF;
    LUT5 ix8473z1315 (.O (nx8473z3), .I0 (\p_sortie_rsc_addr_1_0(0)  ), .I1 (
         \p_rows_rsc_z_int(0)  ), .I2 (\p_fsm_output(8)  ), .I3 (
         \p_fsm_output(0)  ), .I4 (px1473)) ;
         defparam ix8473z1315.INIT = 32'hB3A0FFFF;
endmodule

