mgc_hls.mgc_io_sync_v1(beh) :0:
