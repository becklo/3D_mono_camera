
//------> /softl3/catapultc10_0a/64bit/Mgc_home/pkgs/siflibs/mgc_io_sync_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v1 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


module mgc_in_sync_v1 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0a/269363 Production Release
//  HLS Date:       Wed Nov  9 17:38:00 PST 2016
// 
//  Generated by:   xph3sle509@ocaepc57
//  Generated date: Mon Jan 29 11:55:59 2018
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Xilinx_RAMS_BLOCK_1R1W_RBW_wport_32_17_66880_2_gen
// ------------------------------------------------------------------


module Xilinx_RAMS_BLOCK_1R1W_RBW_wport_32_17_66880_2_gen (
  we, d, wadr, wadr_d, d_d, we_d
);
  output we;
  output [31:0] d;
  output [16:0] wadr;
  input [16:0] wadr_d;
  input [31:0] d_d;
  input we_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_17_66880_1_gen
// ------------------------------------------------------------------


module Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_17_66880_1_gen (
  re, q, radr, radr_d, re_d, q_d
);
  output re;
  input [31:0] q;
  output [16:0] radr;
  input [16:0] radr_d;
  input re_d;
  output [31:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module conv_core_core_fsm (
  clk, rst, fsm_output, for_for_C_2_tr0, for_C_0_tr0
);
  input clk;
  input rst;
  output [5:0] fsm_output;
  reg [5:0] fsm_output;
  input for_for_C_2_tr0;
  input for_C_0_tr0;


  // FSM State Type Declaration for conv_core_core_fsm_1
  parameter
    main_C_0 = 3'd0,
    for_for_C_0 = 3'd1,
    for_for_C_1 = 3'd2,
    for_for_C_2 = 3'd3,
    for_C_0 = 3'd4,
    main_C_1 = 3'd5;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : conv_core_core_fsm_1
    case (state_var)
      for_for_C_0 : begin
        fsm_output = 6'b10;
        state_var_NS = for_for_C_1;
      end
      for_for_C_1 : begin
        fsm_output = 6'b100;
        state_var_NS = for_for_C_2;
      end
      for_for_C_2 : begin
        fsm_output = 6'b1000;
        if ( for_for_C_2_tr0 ) begin
          state_var_NS = for_C_0;
        end
        else begin
          state_var_NS = for_for_C_0;
        end
      end
      for_C_0 : begin
        fsm_output = 6'b10000;
        if ( for_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 6'b100000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 6'b1;
        state_var_NS = for_for_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv_core
// ------------------------------------------------------------------


module conv_core (
  clk, rst, image_in_rsc_triosy_lz, image_out_rsc_triosy_lz, image_in_rsci_radr_d,
      image_in_rsci_re_d, image_in_rsci_q_d, image_out_rsci_wadr_d, image_out_rsci_d_d,
      image_out_rsci_we_d
);
  input clk;
  input rst;
  output image_in_rsc_triosy_lz;
  output image_out_rsc_triosy_lz;
  output [16:0] image_in_rsci_radr_d;
  output image_in_rsci_re_d;
  input [31:0] image_in_rsci_q_d;
  output [16:0] image_out_rsci_wadr_d;
  output [31:0] image_out_rsci_d_d;
  output image_out_rsci_we_d;


  // Interconnect Declarations
  wire [5:0] fsm_output;
  reg [7:0] for_i_7_0_sva_3;
  reg [8:0] for_for_j_8_0_sva_3;
  reg [16:0] for_for_for_for_acc_1_cse_sva;
  reg [8:0] for_for_j_8_0_sva_4;
  reg for_for_slc_for_for_acc_3_itm;
  wire or_2_cse;
  reg reg_image_out_rsc_triosy_obj_ld_cse;
  wire [16:0] for_for_for_for_acc_1_cse_sva_mx0w1;
  wire [17:0] nl_for_for_for_for_acc_1_cse_sva_mx0w1;
  wire [7:0] for_i_7_0_sva_1;
  wire [8:0] nl_for_i_7_0_sva_1;
  wire [8:0] for_for_j_8_0_sva_1;
  wire [9:0] nl_for_for_j_8_0_sva_1;
  wire for_acc_itm_8;

  wire[0:0] not_nl;
  wire[3:0] for_for_acc_nl;
  wire[4:0] nl_for_for_acc_nl;
  wire[16:0] for_for_mul_1_nl;
  wire[8:0] for_acc_nl;
  wire[9:0] nl_for_acc_nl;
  wire[23:0] for_for_for_for_and_nl;
  wire[23:0] for_for_acc_4_nl;
  wire[24:0] nl_for_for_acc_4_nl;
  wire[7:0] for_i_for_i_nor_nl;
  wire[0:0] for_i_not_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_conv_core_core_fsm_inst_for_for_C_2_tr0;
  assign nl_conv_core_core_fsm_inst_for_for_C_2_tr0 = ~ for_for_slc_for_for_acc_3_itm;
  wire [0:0] nl_conv_core_core_fsm_inst_for_C_0_tr0;
  assign nl_conv_core_core_fsm_inst_for_C_0_tr0 = ~ for_acc_itm_8;
  mgc_io_sync_v1 #(.valid(32'sd0)) image_in_rsc_triosy_obj (
      .ld(reg_image_out_rsc_triosy_obj_ld_cse),
      .lz(image_in_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) image_out_rsc_triosy_obj (
      .ld(reg_image_out_rsc_triosy_obj_ld_cse),
      .lz(image_out_rsc_triosy_lz)
    );
  conv_core_core_fsm conv_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .for_for_C_2_tr0(nl_conv_core_core_fsm_inst_for_for_C_2_tr0[0:0]),
      .for_C_0_tr0(nl_conv_core_core_fsm_inst_for_C_0_tr0[0:0])
    );
  assign or_2_cse = (fsm_output[0]) | (fsm_output[4]);
  assign nl_for_i_7_0_sva_1 = for_i_7_0_sva_3 + 8'b1;
  assign for_i_7_0_sva_1 = nl_for_i_7_0_sva_1[7:0];
  assign for_for_mul_1_nl = conv_u2u_17_17((for_for_j_8_0_sva_3) * 8'b11010001);
  assign nl_for_for_for_for_acc_1_cse_sva_mx0w1 = (for_for_mul_1_nl) + conv_u2u_8_17(for_i_7_0_sva_3);
  assign for_for_for_for_acc_1_cse_sva_mx0w1 = nl_for_for_for_for_acc_1_cse_sva_mx0w1[16:0];
  assign nl_for_for_j_8_0_sva_1 = for_for_j_8_0_sva_3 + 9'b1;
  assign for_for_j_8_0_sva_1 = nl_for_for_j_8_0_sva_1[8:0];
  assign nl_for_acc_nl = conv_u2s_8_9(for_i_7_0_sva_1) + 9'b100101111;
  assign for_acc_nl = nl_for_acc_nl[8:0];
  assign for_acc_itm_8 = readslicef_9_1_8((for_acc_nl));
  assign image_in_rsci_radr_d = MUX_v_17_2_2(17'b00000000000000000, for_for_for_for_acc_1_cse_sva_mx0w1,
      (fsm_output[1]));
  assign image_in_rsci_re_d = fsm_output[1];
  assign image_out_rsci_wadr_d = MUX_v_17_2_2(17'b00000000000000000, for_for_for_for_acc_1_cse_sva,
      (fsm_output[2]));
  assign nl_for_for_acc_4_nl =  -(image_in_rsci_q_d[31:8]);
  assign for_for_acc_4_nl = nl_for_for_acc_4_nl[23:0];
  assign for_for_for_for_and_nl = MUX_v_24_2_2(24'b000000000000000000000000, (for_for_acc_4_nl),
      (fsm_output[2]));
  assign for_i_not_nl = ~ (fsm_output[2]);
  assign for_i_for_i_nor_nl = ~(MUX_v_8_2_2((image_in_rsci_q_d[7:0]), 8'b11111111,
      (for_i_not_nl)));
  assign image_out_rsci_d_d = {(for_for_for_for_and_nl) , (for_i_for_i_nor_nl)};
  assign image_out_rsci_we_d = fsm_output[2];
  always @(posedge clk) begin
    if ( rst ) begin
      for_i_7_0_sva_3 <= 8'b0;
    end
    else if ( or_2_cse ) begin
      for_i_7_0_sva_3 <= MUX_v_8_2_2(8'b00000000, for_i_7_0_sva_1, (fsm_output[4]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_j_8_0_sva_3 <= 9'b0;
      reg_image_out_rsc_triosy_obj_ld_cse <= 1'b0;
      for_for_for_for_acc_1_cse_sva <= 17'b0;
    end
    else begin
      for_for_j_8_0_sva_3 <= MUX_v_9_2_2(9'b000000000, for_for_j_8_0_sva_4, (not_nl));
      reg_image_out_rsc_triosy_obj_ld_cse <= (~ for_acc_itm_8) & (fsm_output[4]);
      for_for_for_for_acc_1_cse_sva <= for_for_for_for_acc_1_cse_sva_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_slc_for_for_acc_3_itm <= 1'b0;
    end
    else if ( fsm_output[1] ) begin
      for_for_slc_for_for_acc_3_itm <= readslicef_4_1_3((for_for_acc_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_j_8_0_sva_4 <= 9'b0;
    end
    else if ( fsm_output[1] ) begin
      for_for_j_8_0_sva_4 <= for_for_j_8_0_sva_1;
    end
  end
  assign not_nl = ~ or_2_cse;
  assign nl_for_for_acc_nl = conv_u2s_3_4(for_for_j_8_0_sva_1[8:6]) + 4'b1011;
  assign for_for_acc_nl = nl_for_for_acc_nl[3:0];

  function [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [0:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function  [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function  [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function  [16:0] conv_u2u_8_17 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_17 = {{9{1'b0}}, vector};
  end
  endfunction


  function  [16:0] conv_u2u_17_17 ;
    input [16:0]  vector ;
  begin
    conv_u2u_17_17 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv
// ------------------------------------------------------------------


module conv (
  clk, rst, image_in_rsc_radr, image_in_rsc_q, image_in_rsc_re, image_in_rsc_triosy_lz,
      image_out_rsc_wadr, image_out_rsc_d, image_out_rsc_we, image_out_rsc_triosy_lz
);
  input clk;
  input rst;
  output [16:0] image_in_rsc_radr;
  input [31:0] image_in_rsc_q;
  output image_in_rsc_re;
  output image_in_rsc_triosy_lz;
  output [16:0] image_out_rsc_wadr;
  output [31:0] image_out_rsc_d;
  output image_out_rsc_we;
  output image_out_rsc_triosy_lz;


  // Interconnect Declarations
  wire [16:0] image_in_rsci_radr_d;
  wire image_in_rsci_re_d;
  wire [31:0] image_in_rsci_q_d;
  wire [16:0] image_out_rsci_wadr_d;
  wire [31:0] image_out_rsci_d_d;
  wire image_out_rsci_we_d;


  // Interconnect Declarations for Component Instantiations 
  Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_17_66880_1_gen image_in_rsci (
      .re(image_in_rsc_re),
      .q(image_in_rsc_q),
      .radr(image_in_rsc_radr),
      .radr_d(image_in_rsci_radr_d),
      .re_d(image_in_rsci_re_d),
      .q_d(image_in_rsci_q_d)
    );
  Xilinx_RAMS_BLOCK_1R1W_RBW_wport_32_17_66880_2_gen image_out_rsci (
      .we(image_out_rsc_we),
      .d(image_out_rsc_d),
      .wadr(image_out_rsc_wadr),
      .wadr_d(image_out_rsci_wadr_d),
      .d_d(image_out_rsci_d_d),
      .we_d(image_out_rsci_we_d)
    );
  conv_core conv_core_inst (
      .clk(clk),
      .rst(rst),
      .image_in_rsc_triosy_lz(image_in_rsc_triosy_lz),
      .image_out_rsc_triosy_lz(image_out_rsc_triosy_lz),
      .image_in_rsci_radr_d(image_in_rsci_radr_d),
      .image_in_rsci_re_d(image_in_rsci_re_d),
      .image_in_rsci_q_d(image_in_rsci_q_d),
      .image_out_rsci_wadr_d(image_out_rsci_wadr_d),
      .image_out_rsci_d_d(image_out_rsci_d_d),
      .image_out_rsci_we_d(image_out_rsci_we_d)
    );
endmodule



