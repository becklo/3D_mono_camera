
//------> /softl3/catapultc10_0a/64bit/Mgc_home/pkgs/siflibs/mgc_in_wire_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_wire_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule


//------> /softl3/catapultc10_0a/64bit/Mgc_home/pkgs/siflibs/mgc_io_sync_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v1 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


module mgc_in_sync_v1 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0a/269363 Production Release
//  HLS Date:       Wed Nov  9 17:38:00 PST 2016
// 
//  Generated by:   xph3sle509@ocaepc57
//  Generated date: Tue Jan 23 11:05:31 2018
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rwport_5_68256_32_17_0_1_0_0_0_1_1_1_0_68256_32_1_gen
// ------------------------------------------------------------------


module ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rwport_5_68256_32_17_0_1_0_0_0_1_1_1_0_68256_32_1_gen
    (
  data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d
);
  input [31:0] data_out;
  output we;
  output re;
  output [16:0] addr;
  output [31:0] data_in;
  input [31:0] data_in_d;
  input [16:0] addr_d;
  input re_d;
  input we_d;
  output [31:0] data_out_d;



  // Interconnect Declarations for Component Instantiations 
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rport_4_289_32_9_0_1_0_0_0_1_1_1_0_289_32_1_gen
// ------------------------------------------------------------------


module ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rport_4_289_32_9_0_1_0_0_0_1_1_1_0_289_32_1_gen
    (
  data_out, re, addr, addr_d, re_d, data_out_d
);
  input [31:0] data_out;
  output re;
  output [8:0] addr;
  input [8:0] addr_d;
  input re_d;
  output [31:0] data_out_d;



  // Interconnect Declarations for Component Instantiations 
  assign data_out_d = data_out;
  assign re = (re_d);
  assign addr = (addr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rport_1_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
// ------------------------------------------------------------------


module ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rport_1_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
    (
  data_out, re, addr, addr_d, re_d, data_out_d
);
  input [31:0] data_out;
  output re;
  output [15:0] addr;
  input [15:0] addr_d;
  input re_d;
  output [31:0] data_out_d;



  // Interconnect Declarations for Component Instantiations 
  assign data_out_d = data_out;
  assign re = (re_d);
  assign addr = (addr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module conv_core_core_fsm (
  clk, rst, fsm_output, main_C_0_tr0, for_C_0_tr0, for_for_for_for_C_3_tr0, for_for_for_C_1_tr0,
      for_for_C_0_tr0, for_C_1_tr0
);
  input clk;
  input rst;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;
  input main_C_0_tr0;
  input for_C_0_tr0;
  input for_for_for_for_C_3_tr0;
  input for_for_for_C_1_tr0;
  input for_for_C_0_tr0;
  input for_C_1_tr0;


  // FSM State Type Declaration for conv_core_core_fsm_1
  parameter
    main_C_0 = 4'd0,
    for_C_0 = 4'd1,
    for_for_for_C_0 = 4'd2,
    for_for_for_for_C_0 = 4'd3,
    for_for_for_for_C_1 = 4'd4,
    for_for_for_for_C_2 = 4'd5,
    for_for_for_for_C_3 = 4'd6,
    for_for_for_C_1 = 4'd7,
    for_for_C_0 = 4'd8,
    for_C_1 = 4'd9,
    main_C_1 = 4'd10;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : conv_core_core_fsm_1
    case (state_var)
      for_C_0 : begin
        fsm_output = 11'b10;
        if ( for_C_0_tr0 ) begin
          state_var_NS = for_C_1;
        end
        else begin
          state_var_NS = for_for_for_C_0;
        end
      end
      for_for_for_C_0 : begin
        fsm_output = 11'b100;
        state_var_NS = for_for_for_for_C_0;
      end
      for_for_for_for_C_0 : begin
        fsm_output = 11'b1000;
        state_var_NS = for_for_for_for_C_1;
      end
      for_for_for_for_C_1 : begin
        fsm_output = 11'b10000;
        state_var_NS = for_for_for_for_C_2;
      end
      for_for_for_for_C_2 : begin
        fsm_output = 11'b100000;
        state_var_NS = for_for_for_for_C_3;
      end
      for_for_for_for_C_3 : begin
        fsm_output = 11'b1000000;
        if ( for_for_for_for_C_3_tr0 ) begin
          state_var_NS = for_for_for_C_1;
        end
        else begin
          state_var_NS = for_for_for_for_C_0;
        end
      end
      for_for_for_C_1 : begin
        fsm_output = 11'b10000000;
        if ( for_for_for_C_1_tr0 ) begin
          state_var_NS = for_for_C_0;
        end
        else begin
          state_var_NS = for_for_for_C_0;
        end
      end
      for_for_C_0 : begin
        fsm_output = 11'b100000000;
        if ( for_for_C_0_tr0 ) begin
          state_var_NS = for_C_1;
        end
        else begin
          state_var_NS = for_for_for_C_0;
        end
      end
      for_C_1 : begin
        fsm_output = 11'b1000000000;
        if ( for_C_1_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 11'b10000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 11'b1;
        if ( main_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv_core
// ------------------------------------------------------------------


module conv_core (
  clk, rst, image_rsc_triosy_lz, rows_rsc_z, rows_rsc_triosy_lz, cols_rsc_z, cols_rsc_triosy_lz,
      kernel_rsc_triosy_lz, sortie_rsc_triosy_lz, image_rsci_addr_d, image_rsci_re_d,
      image_rsci_data_out_d, kernel_rsci_addr_d, kernel_rsci_data_out_d, sortie_rsci_data_in_d,
      sortie_rsci_addr_d, sortie_rsci_we_d, sortie_rsci_data_out_d, kernel_rsci_re_d_pff
);
  input clk;
  input rst;
  output image_rsc_triosy_lz;
  input [31:0] rows_rsc_z;
  output rows_rsc_triosy_lz;
  input [31:0] cols_rsc_z;
  output cols_rsc_triosy_lz;
  output kernel_rsc_triosy_lz;
  output sortie_rsc_triosy_lz;
  output [15:0] image_rsci_addr_d;
  output image_rsci_re_d;
  input [31:0] image_rsci_data_out_d;
  output [8:0] kernel_rsci_addr_d;
  wire [9:0] nl_kernel_rsci_addr_d;
  input [31:0] kernel_rsci_data_out_d;
  output [31:0] sortie_rsci_data_in_d;
  output [16:0] sortie_rsci_addr_d;
  output sortie_rsci_we_d;
  input [31:0] sortie_rsci_data_out_d;
  output kernel_rsci_re_d_pff;


  // Interconnect Declarations
  wire [31:0] rows_rsci_d;
  wire [31:0] cols_rsci_d;
  wire [10:0] fsm_output;
  wire [31:0] for_for_for_for_acc_3_tmp;
  wire [32:0] nl_for_for_for_for_acc_3_tmp;
  wire or_tmp_9;
  reg [31:0] rows_1_sva_2;
  reg [31:0] cols_1_sva_1;
  reg [31:0] for_i_sva;
  reg [31:0] for_for_j_sva;
  reg [4:0] for_for_for_m_4_0_sva_4;
  reg [4:0] for_for_for_acc_1_psp_sva;
  wire [5:0] nl_for_for_for_acc_1_psp_sva;
  reg [4:0] for_for_for_for_n_4_0_sva;
  reg [13:0] for_for_for_for_if_acc_psp_sva_1;
  reg [4:0] for_for_for_for_n_4_0_sva_3;
  reg for_for_for_for_if_for_for_for_for_if_and_2_itm;
  reg [31:0] for_for_for_for_if_asn_7_itm_2;
  reg [12:0] for_for_for_for_if_slc_ii_28_0_itm_2;
  reg [12:0] for_for_for_for_if_slc_jj_15_3_itm_2;
  reg [2:0] for_for_for_for_if_slc_jj_2_0_itm_3;
  reg [31:0] for_for_for_for_if_asn_6_itm_2;
  reg for_for_for_for_slc_for_for_for_for_acc_5_itm;
  wire for_for_for_for_aif_acc_tmp_32;
  wire exit_for_sva_mx0;
  wire exit_for_for_sva_mx0;
  wire [31:0] jj_sva;
  wire [32:0] nl_jj_sva;
  reg reg_sortie_rsc_triosy_obj_ld_cse;
  wire or_cse;
  wire [13:0] for_for_for_for_if_acc_psp_sva;
  wire [14:0] nl_for_for_for_for_if_acc_psp_sva;
  wire [32:0] z_out_1;
  wire [32:0] z_out_2;
  wire [33:0] nl_z_out_2;
  wire [31:0] z_out_4;
  wire [63:0] nl_z_out_4;
  wire z_out_4_1;
  wire [4:0] z_out_3_4_0;
  wire [5:0] nl_z_out_3_4_0;

  wire[1:0] for_for_for_for_acc_17_nl;
  wire[2:0] nl_for_for_for_for_acc_17_nl;
  wire[2:0] for_for_for_for_acc_16_nl;
  wire[3:0] nl_for_for_for_for_acc_16_nl;
  wire[32:0] for_for_for_for_aif_acc_nl;
  wire[33:0] nl_for_for_for_for_aif_acc_nl;
  wire[12:0] for_for_for_for_if_acc_3_nl;
  wire[13:0] nl_for_for_for_for_if_acc_3_nl;
  wire[8:0] for_for_for_for_acc_15_nl;
  wire[9:0] nl_for_for_for_for_acc_15_nl;
  wire[1:0] for_for_for_for_acc_18_nl;
  wire[2:0] nl_for_for_for_for_acc_18_nl;
  wire[13:0] sortie_mux_nl;
  wire[33:0] acc_1_nl;
  wire[34:0] nl_acc_1_nl;
  wire[31:0] for_mux1h_4_nl;
  wire[0:0] for_or_3_nl;
  wire[31:0] for_mux1h_5_nl;
  wire[0:0] for_or_5_nl;
  wire[31:0] for_mux1h_6_nl;
  wire[4:0] for_for_for_mux_3_nl;
  wire[31:0] for_for_for_for_if_mux1h_15_nl;
  wire[31:0] for_for_for_for_if_mux1h_16_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_conv_core_core_fsm_inst_for_for_for_for_C_3_tr0;
  assign nl_conv_core_core_fsm_inst_for_for_for_for_C_3_tr0 = ~ for_for_for_for_slc_for_for_for_for_acc_5_itm;
  wire [0:0] nl_conv_core_core_fsm_inst_for_for_for_C_1_tr0;
  assign nl_conv_core_core_fsm_inst_for_for_for_C_1_tr0 = ~ z_out_4_1;
  mgc_in_wire_v1 #(.rscid(32'sd2),
  .width(32'sd32)) rows_rsci (
      .d(rows_rsci_d),
      .z(rows_rsc_z)
    );
  mgc_in_wire_v1 #(.rscid(32'sd3),
  .width(32'sd32)) cols_rsci (
      .d(cols_rsci_d),
      .z(cols_rsc_z)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) image_rsc_triosy_obj (
      .ld(reg_sortie_rsc_triosy_obj_ld_cse),
      .lz(image_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) rows_rsc_triosy_obj (
      .ld(reg_sortie_rsc_triosy_obj_ld_cse),
      .lz(rows_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) cols_rsc_triosy_obj (
      .ld(reg_sortie_rsc_triosy_obj_ld_cse),
      .lz(cols_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) kernel_rsc_triosy_obj (
      .ld(reg_sortie_rsc_triosy_obj_ld_cse),
      .lz(kernel_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) sortie_rsc_triosy_obj (
      .ld(reg_sortie_rsc_triosy_obj_ld_cse),
      .lz(sortie_rsc_triosy_lz)
    );
  conv_core_core_fsm conv_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .main_C_0_tr0(exit_for_sva_mx0),
      .for_C_0_tr0(exit_for_for_sva_mx0),
      .for_for_for_for_C_3_tr0(nl_conv_core_core_fsm_inst_for_for_for_for_C_3_tr0[0:0]),
      .for_for_for_C_1_tr0(nl_conv_core_core_fsm_inst_for_for_for_C_1_tr0[0:0]),
      .for_for_C_0_tr0(exit_for_for_sva_mx0),
      .for_C_1_tr0(exit_for_sva_mx0)
    );
  assign or_cse = (fsm_output[0]) | (fsm_output[9]);
  assign exit_for_sva_mx0 = MUX_s_1_2_2((~ (z_out_2[32])), (~ (z_out_1[32])), fsm_output[9]);
  assign exit_for_for_sva_mx0 = MUX_s_1_2_2((~ (z_out_2[32])), (~ (z_out_1[32])),
      fsm_output[8]);
  assign nl_for_for_for_for_if_acc_psp_sva = (z_out_4[13:0]) + (for_for_j_sva[16:3]);
  assign for_for_for_for_if_acc_psp_sva = nl_for_for_for_for_if_acc_psp_sva[13:0];
  assign nl_for_for_for_for_acc_17_nl = (for_for_for_for_n_4_0_sva[4:3]) + 2'b11;
  assign for_for_for_for_acc_17_nl = nl_for_for_for_for_acc_17_nl[1:0];
  assign nl_jj_sva = conv_s2s_5_32({(for_for_for_for_acc_17_nl) , (for_for_for_for_n_4_0_sva[2:0])})
      + for_for_j_sva;
  assign jj_sva = nl_jj_sva[31:0];
  assign nl_for_for_for_for_acc_16_nl = conv_u2s_2_3(for_for_for_m_4_0_sva_4[4:3])
      + 3'b111;
  assign for_for_for_for_acc_16_nl = nl_for_for_for_for_acc_16_nl[2:0];
  assign nl_for_for_for_for_acc_3_tmp = conv_s2s_6_32({(for_for_for_for_acc_16_nl)
      , (for_for_for_m_4_0_sva_4[2:0])}) + for_i_sva;
  assign for_for_for_for_acc_3_tmp = nl_for_for_for_for_acc_3_tmp[31:0];
  assign nl_for_for_for_for_aif_acc_nl = conv_u2u_31_33(for_for_for_for_acc_3_tmp[30:0])
      - conv_s2u_32_33(rows_1_sva_2);
  assign for_for_for_for_aif_acc_nl = nl_for_for_for_for_aif_acc_nl[32:0];
  assign for_for_for_for_aif_acc_tmp_32 = readslicef_33_1_32((for_for_for_for_aif_acc_nl));
  assign or_tmp_9 = ~((fsm_output[10]) | (fsm_output[0]));
  assign nl_for_for_for_for_if_acc_3_nl = (z_out_4[12:0]) + for_for_for_for_if_slc_jj_15_3_itm_2;
  assign for_for_for_for_if_acc_3_nl = nl_for_for_for_for_if_acc_3_nl[12:0];
  assign image_rsci_addr_d = {(for_for_for_for_if_acc_3_nl) , for_for_for_for_if_slc_jj_2_0_itm_3};
  assign image_rsci_re_d = ~(for_for_for_for_if_for_for_for_for_if_and_2_itm & (fsm_output[4]));
  assign nl_for_for_for_for_acc_18_nl = conv_u2u_1_2(for_for_for_acc_1_psp_sva[4])
      + 2'b1;
  assign for_for_for_for_acc_18_nl = nl_for_for_for_for_acc_18_nl[1:0];
  assign nl_for_for_for_for_acc_15_nl = ({for_for_for_acc_1_psp_sva , 4'b1}) + conv_u2u_6_9({(for_for_for_for_acc_18_nl)
      , (for_for_for_acc_1_psp_sva[3:0])});
  assign for_for_for_for_acc_15_nl = nl_for_for_for_for_acc_15_nl[8:0];
  assign nl_kernel_rsci_addr_d = (for_for_for_for_acc_15_nl) + ({4'b1111 , (~ for_for_for_for_n_4_0_sva)});
  assign kernel_rsci_addr_d = nl_kernel_rsci_addr_d[8:0];
  assign kernel_rsci_re_d_pff = ~((~ (for_for_for_for_acc_3_tmp[31])) & for_for_for_for_aif_acc_tmp_32
      & (~ (jj_sva[31])) & (z_out_1[32]) & (fsm_output[3]));
  assign sortie_mux_nl = MUX_v_14_2_2(for_for_for_for_if_acc_psp_sva, for_for_for_for_if_acc_psp_sva_1,
      fsm_output[5]);
  assign sortie_rsci_addr_d = {(sortie_mux_nl) , (for_for_j_sva[2:0])};
  assign sortie_rsci_we_d = ~(for_for_for_for_if_for_for_for_for_if_and_2_itm & (fsm_output[5]));
  assign sortie_rsci_data_in_d = z_out_1[31:0];
  always @(posedge clk) begin
    if ( rst ) begin
      reg_sortie_rsc_triosy_obj_ld_cse <= 1'b0;
      for_for_for_for_n_4_0_sva <= 5'b0;
      for_for_for_for_if_slc_jj_2_0_itm_3 <= 3'b0;
      for_for_for_for_if_slc_jj_15_3_itm_2 <= 13'b0;
      for_for_for_for_if_slc_ii_28_0_itm_2 <= 13'b0;
      for_for_for_for_if_asn_6_itm_2 <= 32'b0;
      for_for_for_for_if_asn_7_itm_2 <= 32'b0;
    end
    else begin
      reg_sortie_rsc_triosy_obj_ld_cse <= or_cse & exit_for_sva_mx0;
      for_for_for_for_n_4_0_sva <= MUX_v_5_2_2(5'b00000, for_for_for_for_n_4_0_sva_3,
          (fsm_output[6]));
      for_for_for_for_if_slc_jj_2_0_itm_3 <= jj_sva[2:0];
      for_for_for_for_if_slc_jj_15_3_itm_2 <= jj_sva[15:3];
      for_for_for_for_if_slc_ii_28_0_itm_2 <= for_for_for_for_acc_3_tmp[12:0];
      for_for_for_for_if_asn_6_itm_2 <= kernel_rsci_data_out_d;
      for_for_for_for_if_asn_7_itm_2 <= sortie_rsci_data_out_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      rows_1_sva_2 <= 32'b0;
    end
    else if ( ~ or_tmp_9 ) begin
      rows_1_sva_2 <= rows_rsci_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_i_sva <= 32'b0;
    end
    else if ( or_cse ) begin
      for_i_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000, (z_out_2[31:0]),
          (fsm_output[9]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      cols_1_sva_1 <= 32'b0;
    end
    else if ( ~ or_tmp_9 ) begin
      cols_1_sva_1 <= cols_rsci_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_j_sva <= 32'b0;
    end
    else if ( (fsm_output[1]) | (fsm_output[8]) ) begin
      for_for_j_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000, (z_out_2[31:0]),
          (fsm_output[8]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_m_4_0_sva_4 <= 5'b0;
    end
    else if ( (fsm_output[8]) | (fsm_output[1]) | (fsm_output[7]) ) begin
      for_for_for_m_4_0_sva_4 <= MUX_v_5_2_2(5'b00000, z_out_3_4_0, (fsm_output[7]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_acc_1_psp_sva <= 5'b0;
    end
    else if ( ~((fsm_output[6:3]!=4'b0000)) ) begin
      for_for_for_acc_1_psp_sva <= nl_for_for_for_acc_1_psp_sva[4:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_for_if_acc_psp_sva_1 <= 14'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      for_for_for_for_if_acc_psp_sva_1 <= for_for_for_for_if_acc_psp_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_for_slc_for_for_for_for_acc_5_itm <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      for_for_for_for_slc_for_for_for_for_acc_5_itm <= z_out_4_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_for_if_for_for_for_for_if_and_2_itm <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      for_for_for_for_if_for_for_for_for_if_and_2_itm <= (z_out_1[32]) & (~ (jj_sva[31]))
          & for_for_for_for_aif_acc_tmp_32 & (~ (for_for_for_for_acc_3_tmp[31]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_for_n_4_0_sva_3 <= 5'b0;
    end
    else if ( fsm_output[3] ) begin
      for_for_for_for_n_4_0_sva_3 <= z_out_3_4_0;
    end
  end
  assign nl_for_for_for_acc_1_psp_sva  = (~ for_for_for_m_4_0_sva_4) + 5'b10001;
  assign z_out_4_1 = (z_out_3_4_0[4]) ^ ((z_out_3_4_0[3:0]!=4'b0000));
  assign for_or_3_nl = (fsm_output[9:8]!=2'b00);
  assign for_mux1h_4_nl = MUX1HOT_v_32_3_2((z_out_2[31:0]), jj_sva, for_for_for_for_if_asn_7_itm_2,
      {(for_or_3_nl) , (fsm_output[3]) , (fsm_output[5])});
  assign for_or_5_nl = (fsm_output[8]) | (fsm_output[3]);
  assign for_mux1h_5_nl = MUX1HOT_v_32_3_2((~ rows_1_sva_2), (~ cols_1_sva_1), z_out_4,
      {(fsm_output[9]) , (for_or_5_nl) , (fsm_output[5])});
  assign nl_acc_1_nl = conv_s2u_33_34({(for_mux1h_4_nl) , (~ (fsm_output[5]))}) +
      conv_s2u_33_34({(for_mux1h_5_nl) , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[33:0];
  assign z_out_1 = readslicef_34_33_1((acc_1_nl));
  assign for_mux1h_6_nl = MUX1HOT_v_32_4_2((~ rows_rsci_d), for_i_sva, (~ cols_1_sva_1),
      for_for_j_sva, {(fsm_output[0]) , (fsm_output[9]) , (fsm_output[1]) , (fsm_output[8])});
  assign nl_z_out_2 = conv_s2u_32_33(for_mux1h_6_nl) + 33'b1;
  assign z_out_2 = nl_z_out_2[32:0];
  assign for_for_for_mux_3_nl = MUX_v_5_2_2(for_for_for_m_4_0_sva_4, for_for_for_for_n_4_0_sva,
      fsm_output[3]);
  assign nl_z_out_3_4_0 = (for_for_for_mux_3_nl) + 5'b1;
  assign z_out_3_4_0 = nl_z_out_3_4_0[4:0];
  assign for_for_for_for_if_mux1h_15_nl = MUX1HOT_v_32_3_2((signext_32_14(for_i_sva[13:0])),
      ({19'b0 , for_for_for_for_if_slc_ii_28_0_itm_2}), image_rsci_data_out_d, {(fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5])});
  assign for_for_for_for_if_mux1h_16_nl = MUX1HOT_v_32_3_2(32'b11011, 32'b11001,
      for_for_for_for_if_asn_6_itm_2, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_z_out_4 = (for_for_for_for_if_mux1h_15_nl) * (for_for_for_for_if_mux1h_16_nl);
  assign z_out_4 = nl_z_out_4[31:0];

  function [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function [31:0] MUX1HOT_v_32_4_2;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [3:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    MUX1HOT_v_32_4_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function [32:0] readslicef_34_33_1;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_34_33_1 = tmp[32:0];
  end
  endfunction


  function [31:0] signext_32_14;
    input [13:0] vector;
  begin
    signext_32_14= {{18{vector[13]}}, vector};
  end
  endfunction


  function  [31:0] conv_s2s_5_32 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_32 = {{27{vector[4]}}, vector};
  end
  endfunction


  function  [31:0] conv_s2s_6_32 ;
    input [5:0]  vector ;
  begin
    conv_s2s_6_32 = {{26{vector[5]}}, vector};
  end
  endfunction


  function  [32:0] conv_s2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_s2u_32_33 = {vector[31], vector};
  end
  endfunction


  function  [33:0] conv_s2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_s2u_33_34 = {vector[32], vector};
  end
  endfunction


  function  [2:0] conv_u2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2s_2_3 =  {1'b0, vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function  [8:0] conv_u2u_6_9 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_9 = {{3{1'b0}}, vector};
  end
  endfunction


  function  [32:0] conv_u2u_31_33 ;
    input [30:0]  vector ;
  begin
    conv_u2u_31_33 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv
// ------------------------------------------------------------------


module conv (
  clk, rst, image_rsc_addr, image_rsc_re, image_rsc_data_out, image_rsc_triosy_lz,
      rows_rsc_z, rows_rsc_triosy_lz, cols_rsc_z, cols_rsc_triosy_lz, kernel_rsc_addr,
      kernel_rsc_re, kernel_rsc_data_out, kernel_rsc_triosy_lz, sortie_rsc_data_in,
      sortie_rsc_addr, sortie_rsc_re, sortie_rsc_we, sortie_rsc_data_out, sortie_rsc_triosy_lz
);
  input clk;
  input rst;
  output [15:0] image_rsc_addr;
  output image_rsc_re;
  input [31:0] image_rsc_data_out;
  output image_rsc_triosy_lz;
  input [31:0] rows_rsc_z;
  output rows_rsc_triosy_lz;
  input [31:0] cols_rsc_z;
  output cols_rsc_triosy_lz;
  output [8:0] kernel_rsc_addr;
  output kernel_rsc_re;
  input [31:0] kernel_rsc_data_out;
  output kernel_rsc_triosy_lz;
  output [31:0] sortie_rsc_data_in;
  output [16:0] sortie_rsc_addr;
  output sortie_rsc_re;
  output sortie_rsc_we;
  input [31:0] sortie_rsc_data_out;
  output sortie_rsc_triosy_lz;


  // Interconnect Declarations
  wire [15:0] image_rsci_addr_d;
  wire image_rsci_re_d;
  wire [31:0] image_rsci_data_out_d;
  wire [8:0] kernel_rsci_addr_d;
  wire [31:0] kernel_rsci_data_out_d;
  wire [31:0] sortie_rsci_data_in_d;
  wire [16:0] sortie_rsci_addr_d;
  wire sortie_rsci_we_d;
  wire [31:0] sortie_rsci_data_out_d;
  wire kernel_rsci_re_d_iff;


  // Interconnect Declarations for Component Instantiations 
  ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rport_1_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
      image_rsci (
      .data_out(image_rsc_data_out),
      .re(image_rsc_re),
      .addr(image_rsc_addr),
      .addr_d(image_rsci_addr_d),
      .re_d(image_rsci_re_d),
      .data_out_d(image_rsci_data_out_d)
    );
  ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rport_4_289_32_9_0_1_0_0_0_1_1_1_0_289_32_1_gen
      kernel_rsci (
      .data_out(kernel_rsc_data_out),
      .re(kernel_rsc_re),
      .addr(kernel_rsc_addr),
      .addr_d(kernel_rsci_addr_d),
      .re_d(kernel_rsci_re_d_iff),
      .data_out_d(kernel_rsci_data_out_d)
    );
  ram_Xilinx_ARTIX_7_3_RAMSB_singleport_rwport_5_68256_32_17_0_1_0_0_0_1_1_1_0_68256_32_1_gen
      sortie_rsci (
      .data_out(sortie_rsc_data_out),
      .we(sortie_rsc_we),
      .re(sortie_rsc_re),
      .addr(sortie_rsc_addr),
      .data_in(sortie_rsc_data_in),
      .data_in_d(sortie_rsci_data_in_d),
      .addr_d(sortie_rsci_addr_d),
      .re_d(kernel_rsci_re_d_iff),
      .we_d(sortie_rsci_we_d),
      .data_out_d(sortie_rsci_data_out_d)
    );
  conv_core conv_core_inst (
      .clk(clk),
      .rst(rst),
      .image_rsc_triosy_lz(image_rsc_triosy_lz),
      .rows_rsc_z(rows_rsc_z),
      .rows_rsc_triosy_lz(rows_rsc_triosy_lz),
      .cols_rsc_z(cols_rsc_z),
      .cols_rsc_triosy_lz(cols_rsc_triosy_lz),
      .kernel_rsc_triosy_lz(kernel_rsc_triosy_lz),
      .sortie_rsc_triosy_lz(sortie_rsc_triosy_lz),
      .image_rsci_addr_d(image_rsci_addr_d),
      .image_rsci_re_d(image_rsci_re_d),
      .image_rsci_data_out_d(image_rsci_data_out_d),
      .kernel_rsci_addr_d(kernel_rsci_addr_d),
      .kernel_rsci_data_out_d(kernel_rsci_data_out_d),
      .sortie_rsci_data_in_d(sortie_rsci_data_in_d),
      .sortie_rsci_addr_d(sortie_rsci_addr_d),
      .sortie_rsci_we_d(sortie_rsci_we_d),
      .sortie_rsci_data_out_d(sortie_rsci_data_out_d),
      .kernel_rsci_re_d_pff(kernel_rsci_re_d_iff)
    );
endmodule



