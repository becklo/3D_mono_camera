
//------> /softl3/catapultc10_0a/64bit/Mgc_home/pkgs/siflibs/mgc_out_stdreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module mgc_out_stdreg_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule




//------> /softl3/catapultc10_0a/64bit/Mgc_home/pkgs/siflibs/mgc_io_sync_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v1 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


module mgc_in_sync_v1 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0a/269363 Production Release
//  HLS Date:       Wed Nov  9 17:38:00 PST 2016
// 
//  Generated by:   xph3sle509@ocaepc57
//  Generated date: Tue Jan 16 14:33:19 2018
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ram_Xilinx_KINTEX_7_3_RAMSB_singleport_wport_6_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
// ------------------------------------------------------------------


module ram_Xilinx_KINTEX_7_3_RAMSB_singleport_wport_6_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
    (
  we, addr, data_in, data_in_d, addr_d, we_d
);
  output we;
  output [15:0] addr;
  output [31:0] data_in;
  input [31:0] data_in_d;
  input [15:0] addr_d;
  input we_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rwport_5_68256_32_17_0_1_0_0_0_1_1_1_0_68256_32_1_gen
// ------------------------------------------------------------------


module ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rwport_5_68256_32_17_0_1_0_0_0_1_1_1_0_68256_32_1_gen
    (
  data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d
);
  input [31:0] data_out;
  output we;
  output re;
  output [16:0] addr;
  output [31:0] data_in;
  input [31:0] data_in_d;
  input [16:0] addr_d;
  input re_d;
  input we_d;
  output [31:0] data_out_d;



  // Interconnect Declarations for Component Instantiations 
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rport_4_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
// ------------------------------------------------------------------


module ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rport_4_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
    (
  data_out, re, addr, addr_d, re_d, data_out_d
);
  input [31:0] data_out;
  output re;
  output [15:0] addr;
  input [15:0] addr_d;
  input re_d;
  output [31:0] data_out_d;



  // Interconnect Declarations for Component Instantiations 
  assign data_out_d = data_out;
  assign re = (re_d);
  assign addr = (addr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rport_3_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
// ------------------------------------------------------------------


module ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rport_3_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
    (
  data_out, re, addr, addr_d, re_d, data_out_d
);
  input [31:0] data_out;
  output re;
  output [15:0] addr;
  input [15:0] addr_d;
  input re_d;
  output [31:0] data_out_d;



  // Interconnect Declarations for Component Instantiations 
  assign data_out_d = data_out;
  assign re = (re_d);
  assign addr = (addr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    main_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module main_core_core_fsm (
  clk, rst, fsm_output, for_for_C_2_tr0, for_C_0_tr0, for_1_for_C_0_tr0, reconstruction_error_for_C_0_tr0,
      reconstruction_error_for_for_C_1_tr0, reconstruction_error_for_C_1_tr0, for_1_for_C_2_tr0,
      for_1_C_0_tr0
);
  input clk;
  input rst;
  output [13:0] fsm_output;
  reg [13:0] fsm_output;
  input for_for_C_2_tr0;
  input for_C_0_tr0;
  input for_1_for_C_0_tr0;
  input reconstruction_error_for_C_0_tr0;
  input reconstruction_error_for_for_C_1_tr0;
  input reconstruction_error_for_C_1_tr0;
  input for_1_for_C_2_tr0;
  input for_1_C_0_tr0;


  // FSM State Type Declaration for main_core_core_fsm_1
  parameter
    main_C_0 = 4'd0,
    for_for_C_0 = 4'd1,
    for_for_C_1 = 4'd2,
    for_for_C_2 = 4'd3,
    for_C_0 = 4'd4,
    for_1_for_C_0 = 4'd5,
    reconstruction_error_for_C_0 = 4'd6,
    reconstruction_error_for_for_C_0 = 4'd7,
    reconstruction_error_for_for_C_1 = 4'd8,
    reconstruction_error_for_C_1 = 4'd9,
    for_1_for_C_1 = 4'd10,
    for_1_for_C_2 = 4'd11,
    for_1_C_0 = 4'd12,
    main_C_1 = 4'd13;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : main_core_core_fsm_1
    case (state_var)
      for_for_C_0 : begin
        fsm_output = 14'b10;
        state_var_NS = for_for_C_1;
      end
      for_for_C_1 : begin
        fsm_output = 14'b100;
        state_var_NS = for_for_C_2;
      end
      for_for_C_2 : begin
        fsm_output = 14'b1000;
        if ( for_for_C_2_tr0 ) begin
          state_var_NS = for_C_0;
        end
        else begin
          state_var_NS = for_for_C_0;
        end
      end
      for_C_0 : begin
        fsm_output = 14'b10000;
        if ( for_C_0_tr0 ) begin
          state_var_NS = for_1_for_C_0;
        end
        else begin
          state_var_NS = for_for_C_0;
        end
      end
      for_1_for_C_0 : begin
        fsm_output = 14'b100000;
        if ( for_1_for_C_0_tr0 ) begin
          state_var_NS = for_1_for_C_1;
        end
        else begin
          state_var_NS = reconstruction_error_for_C_0;
        end
      end
      reconstruction_error_for_C_0 : begin
        fsm_output = 14'b1000000;
        if ( reconstruction_error_for_C_0_tr0 ) begin
          state_var_NS = reconstruction_error_for_C_1;
        end
        else begin
          state_var_NS = reconstruction_error_for_for_C_0;
        end
      end
      reconstruction_error_for_for_C_0 : begin
        fsm_output = 14'b10000000;
        state_var_NS = reconstruction_error_for_for_C_1;
      end
      reconstruction_error_for_for_C_1 : begin
        fsm_output = 14'b100000000;
        if ( reconstruction_error_for_for_C_1_tr0 ) begin
          state_var_NS = reconstruction_error_for_C_1;
        end
        else begin
          state_var_NS = reconstruction_error_for_for_C_0;
        end
      end
      reconstruction_error_for_C_1 : begin
        fsm_output = 14'b1000000000;
        if ( reconstruction_error_for_C_1_tr0 ) begin
          state_var_NS = for_1_for_C_1;
        end
        else begin
          state_var_NS = reconstruction_error_for_C_0;
        end
      end
      for_1_for_C_1 : begin
        fsm_output = 14'b10000000000;
        state_var_NS = for_1_for_C_2;
      end
      for_1_for_C_2 : begin
        fsm_output = 14'b100000000000;
        if ( for_1_for_C_2_tr0 ) begin
          state_var_NS = for_1_C_0;
        end
        else begin
          state_var_NS = for_1_for_C_0;
        end
      end
      for_1_C_0 : begin
        fsm_output = 14'b1000000000000;
        if ( for_1_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_1_for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 14'b10000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 14'b1;
        state_var_NS = for_for_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    main_core
// ------------------------------------------------------------------


module main_core (
  clk, rst, image_net_rsc_triosy_lz, image_floue_rsc_triosy_lz, image_error_rsc_triosy_lz,
      depth_rsc_triosy_lz, return_rsc_z, return_rsc_triosy_lz, image_net_rsci_addr_d,
      image_net_rsci_data_out_d, image_floue_rsci_addr_d, image_floue_rsci_data_out_d,
      image_error_rsci_data_in_d, image_error_rsci_addr_d, image_error_rsci_re_d,
      image_error_rsci_we_d, image_error_rsci_data_out_d, depth_rsci_data_in_d, depth_rsci_addr_d,
      depth_rsci_we_d, image_net_rsci_re_d_pff
);
  input clk;
  input rst;
  output image_net_rsc_triosy_lz;
  output image_floue_rsc_triosy_lz;
  output image_error_rsc_triosy_lz;
  output depth_rsc_triosy_lz;
  output [31:0] return_rsc_z;
  output return_rsc_triosy_lz;
  output [15:0] image_net_rsci_addr_d;
  input [31:0] image_net_rsci_data_out_d;
  output [15:0] image_floue_rsci_addr_d;
  input [31:0] image_floue_rsci_data_out_d;
  output [31:0] image_error_rsci_data_in_d;
  output [16:0] image_error_rsci_addr_d;
  output image_error_rsci_re_d;
  output image_error_rsci_we_d;
  input [31:0] image_error_rsci_data_out_d;
  output [31:0] depth_rsci_data_in_d;
  output [15:0] depth_rsci_addr_d;
  output depth_rsci_we_d;
  output image_net_rsci_re_d_pff;


  // Interconnect Declarations
  wire [13:0] fsm_output;
  wire or_tmp_30;
  reg [7:0] for_i_7_0_sva_3;
  reg [8:0] for_for_j_8_0_sva_3;
  reg [8:0] for_for_j_8_0_sva_4;
  reg [7:0] for_1_i_7_0_sva_4;
  reg [8:0] for_1_for_j_8_0_sva;
  reg [4:0] for_1_for_acc_6_psp_1_sva_1;
  reg [5:0] for_1_for_acc_7_psp_1_sva_1;
  wire [6:0] nl_for_1_for_acc_7_psp_1_sva_1;
  reg [31:0] reconstruction_error_rec_error_sva;
  reg [31:0] reconstruction_error_for_l_sva_3;
  reg [31:0] reconstruction_error_rec_error_lpi_6;
  reg exit_reconstruction_error_for_for_sva_1;
  reg [8:0] for_1_for_j_8_0_sva_4;
  reg for_for_if_for_for_if_and_itm_1;
  reg [13:0] for_for_else_acc_itm_2;
  wire [14:0] nl_for_for_else_acc_itm_2;
  reg for_for_slc_for_for_acc_7_itm;
  reg for_1_for_slc_for_1_for_acc_7_itm_1;
  reg [22:0] reconstruction_error_for_for_c_sva_31_9_2;
  reg [8:0] reconstruction_error_for_for_c_sva_8_0_2;
  wire for_for_if_acc_1_tmp_5;
  wire exit_reconstruction_error_for_sva_mx0;
  wire [13:0] reconstruction_error_for_for_acc_6_sdt;
  wire [14:0] nl_reconstruction_error_for_for_acc_6_sdt;
  reg reg_return_rsc_triosy_obj_ld_cse;
  wire or_11_cse;
  wire or_10_cse;
  wire or_18_cse;
  wire [31:0] z_out;
  wire [63:0] nl_z_out;
  wire [12:0] z_out_1;
  wire [13:0] nl_z_out_1;
  wire [7:0] z_out_2;
  wire [8:0] nl_z_out_2;
  wire [7:0] z_out_3;
  wire [8:0] nl_z_out_3;
  wire [6:0] z_out_4;
  wire [7:0] nl_z_out_4;
  wire [8:0] z_out_5;
  wire [9:0] nl_z_out_5;
  wire [31:0] z_out_6;
  wire [31:0] z_out_8;
  wire [32:0] nl_z_out_8;
  wire [4:0] for_1_for_acc_6_psp_1_sva;
  wire [5:0] nl_for_1_for_acc_6_psp_1_sva;
  wire [7:0] reconstruction_error_for_l_acc_psp;
  wire [8:0] nl_reconstruction_error_for_l_acc_psp;
  wire [8:0] reconstruction_error_for_for_c_acc_psp;
  wire [9:0] nl_reconstruction_error_for_for_c_acc_psp;
  wire for_for_aif_oif_acc_itm_9;
  wire for_for_oif_acc_itm_8;
  wire z_out_7_32;
  wire z_out_9_5;

  wire[0:0] not_39_nl;
  wire[31:0] reconstruction_error_rec_error_mux1h_4_nl;
  wire[0:0] not_34_nl;
  wire[31:0] reconstruction_error_rec_error_mux1h_5_nl;
  wire[0:0] or_49_nl;
  wire[0:0] not_nl;
  wire[22:0] reconstruction_error_for_for_c_mux_nl;
  wire[0:0] not_38_nl;
  wire[9:0] for_for_aif_oif_acc_nl;
  wire[10:0] nl_for_for_aif_oif_acc_nl;
  wire[8:0] for_for_oif_acc_nl;
  wire[9:0] nl_for_for_oif_acc_nl;
  wire[5:0] for_for_if_acc_1_nl;
  wire[6:0] nl_for_for_if_acc_1_nl;
  wire[8:0] reconstruction_error_for_acc_3_nl;
  wire[9:0] nl_reconstruction_error_for_acc_3_nl;
  wire[0:0] image_error_mux1h_nl;
  wire[3:0] image_error_image_error_and_nl;
  wire[3:0] image_error_mux_nl;
  wire[0:0] image_error_not_2_nl;
  wire[8:0] image_error_mux1h_2_nl;
  wire[8:0] for_for_if_acc_nl;
  wire[9:0] nl_for_for_if_acc_nl;
  wire[2:0] image_error_image_error_mux_nl;
  wire[17:0] reconstruction_error_for_for_reconstruction_error_for_for_and_2_nl;
  wire[0:0] reconstruction_error_for_for_nor_2_nl;
  wire[4:0] reconstruction_error_for_for_reconstruction_error_for_for_and_3_nl;
  wire[4:0] reconstruction_error_for_for_mux_3_nl;
  wire[0:0] reconstruction_error_for_for_nor_3_nl;
  wire[8:0] reconstruction_error_for_for_mux1h_2_nl;
  wire[31:0] reconstruction_error_for_for_mux1h_3_nl;
  wire[0:0] reconstruction_error_for_for_or_2_nl;
  wire[12:0] for_for_else_mux_2_nl;
  wire[12:0] for_for_else_mul_2_nl;
  wire[13:0] nl_for_for_else_mul_2_nl;
  wire[4:0] for_for_else_mux_3_nl;
  wire[7:0] for_for_mux1h_2_nl;
  wire[6:0] mux_2_nl;
  wire[0:0] or_60_nl;
  wire[7:0] for_mux_3_nl;
  wire[5:0] for_for_aelse_mux_4_nl;
  wire[8:0] for_for_mux_2_nl;
  wire[32:0] acc_5_nl;
  wire[33:0] nl_acc_5_nl;
  wire[31:0] reconstruction_error_for_for_mux_4_nl;
  wire[31:0] reconstruction_error_for_for_mux_5_nl;
  wire[32:0] reconstruction_error_for_acc_nl;
  wire[33:0] nl_reconstruction_error_for_acc_nl;
  wire[31:0] reconstruction_error_for_reconstruction_error_for_mux_1_nl;
  wire[0:0] reconstruction_error_for_reconstruction_error_for_or_1_nl;
  wire[5:0] reconstruction_error_for_reconstruction_error_for_and_1_nl;
  wire[5:0] reconstruction_error_for_mux_4_nl;
  wire[5:0] reconstruction_error_for_acc_8_nl;
  wire[6:0] nl_reconstruction_error_for_acc_8_nl;
  wire[0:0] reconstruction_error_for_not_13_nl;
  wire[1:0] reconstruction_error_for_mux1h_2_nl;
  wire[31:0] reconstruction_error_for_mux_5_nl;
  wire[5:0] for_acc_nl;
  wire[6:0] nl_for_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_main_core_core_fsm_inst_for_for_C_2_tr0;
  assign nl_main_core_core_fsm_inst_for_for_C_2_tr0 = ~ for_for_slc_for_for_acc_7_itm;
  wire [0:0] nl_main_core_core_fsm_inst_for_C_0_tr0;
  assign nl_main_core_core_fsm_inst_for_C_0_tr0 = ~ z_out_9_5;
  wire[7:0] reconstruction_error_for_for_acc_10_nl;
  wire[8:0] nl_reconstruction_error_for_for_acc_10_nl;
  wire[9:0] reconstruction_error_for_for_acc_8_nl;
  wire[10:0] nl_reconstruction_error_for_for_acc_8_nl;
  wire [0:0] nl_main_core_core_fsm_inst_reconstruction_error_for_C_0_tr0;
  assign nl_reconstruction_error_for_for_acc_8_nl = conv_u2u_9_10({(~ for_1_for_acc_7_psp_1_sva_1)
      , (~ (for_1_for_j_8_0_sva[2:0]))}) + conv_u2u_9_10(reconstruction_error_for_for_c_acc_psp);
  assign reconstruction_error_for_for_acc_8_nl = nl_reconstruction_error_for_for_acc_8_nl[9:0];
  assign nl_reconstruction_error_for_for_acc_10_nl = (readslicef_10_8_2((reconstruction_error_for_for_acc_8_nl)))
      + 8'b1111111;
  assign reconstruction_error_for_for_acc_10_nl = nl_reconstruction_error_for_for_acc_10_nl[7:0];
  assign nl_main_core_core_fsm_inst_reconstruction_error_for_C_0_tr0 = ~ (readslicef_8_1_7((reconstruction_error_for_for_acc_10_nl)));
  wire [0:0] nl_main_core_core_fsm_inst_for_1_for_C_2_tr0;
  assign nl_main_core_core_fsm_inst_for_1_for_C_2_tr0 = ~ for_1_for_slc_for_1_for_acc_7_itm_1;
  wire [0:0] nl_main_core_core_fsm_inst_for_1_C_0_tr0;
  assign nl_main_core_core_fsm_inst_for_1_C_0_tr0 = ~ z_out_9_5;
  mgc_out_stdreg_v1 #(.rscid(32'sd7),
  .width(32'sd32)) return_rsci (
      .d(32'b0),
      .z(return_rsc_z)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) image_net_rsc_triosy_obj (
      .ld(reg_return_rsc_triosy_obj_ld_cse),
      .lz(image_net_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) image_floue_rsc_triosy_obj (
      .ld(reg_return_rsc_triosy_obj_ld_cse),
      .lz(image_floue_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) image_error_rsc_triosy_obj (
      .ld(reg_return_rsc_triosy_obj_ld_cse),
      .lz(image_error_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) depth_rsc_triosy_obj (
      .ld(reg_return_rsc_triosy_obj_ld_cse),
      .lz(depth_rsc_triosy_lz)
    );
  mgc_io_sync_v1 #(.valid(32'sd0)) return_rsc_triosy_obj (
      .ld(reg_return_rsc_triosy_obj_ld_cse),
      .lz(return_rsc_triosy_lz)
    );
  main_core_core_fsm main_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .for_for_C_2_tr0(nl_main_core_core_fsm_inst_for_for_C_2_tr0[0:0]),
      .for_C_0_tr0(nl_main_core_core_fsm_inst_for_C_0_tr0[0:0]),
      .for_1_for_C_0_tr0(exit_reconstruction_error_for_sva_mx0),
      .reconstruction_error_for_C_0_tr0(nl_main_core_core_fsm_inst_reconstruction_error_for_C_0_tr0[0:0]),
      .reconstruction_error_for_for_C_1_tr0(exit_reconstruction_error_for_for_sva_1),
      .reconstruction_error_for_C_1_tr0(exit_reconstruction_error_for_sva_mx0),
      .for_1_for_C_2_tr0(nl_main_core_core_fsm_inst_for_1_for_C_2_tr0[0:0]),
      .for_1_C_0_tr0(nl_main_core_core_fsm_inst_for_1_C_0_tr0[0:0])
    );
  assign or_18_cse = (fsm_output[0]) | (fsm_output[4]);
  assign or_11_cse = (z_out_4[6]) | for_for_aif_oif_acc_itm_9;
  assign or_10_cse = for_for_if_acc_1_tmp_5 | for_for_oif_acc_itm_8;
  assign nl_reconstruction_error_for_for_acc_6_sdt = (z_out[13:0]) + (reconstruction_error_for_l_sva_3[16:3]);
  assign reconstruction_error_for_for_acc_6_sdt = nl_reconstruction_error_for_for_acc_6_sdt[13:0];
  assign nl_for_for_aif_oif_acc_nl = ({1'b1 , (~ for_for_j_8_0_sva_3)}) + 10'b100110101;
  assign for_for_aif_oif_acc_nl = nl_for_for_aif_oif_acc_nl[9:0];
  assign for_for_aif_oif_acc_itm_9 = readslicef_10_1_9((for_for_aif_oif_acc_nl));
  assign nl_for_for_oif_acc_nl = ({1'b1 , (~ for_i_7_0_sva_3)}) + 9'b11010001;
  assign for_for_oif_acc_nl = nl_for_for_oif_acc_nl[8:0];
  assign for_for_oif_acc_itm_8 = readslicef_9_1_8((for_for_oif_acc_nl));
  assign nl_for_for_if_acc_1_nl = conv_u2s_5_6(for_i_7_0_sva_3[7:3]) + 6'b111111;
  assign for_for_if_acc_1_nl = nl_for_for_if_acc_1_nl[5:0];
  assign for_for_if_acc_1_tmp_5 = readslicef_6_1_5((for_for_if_acc_1_nl));
  assign nl_reconstruction_error_for_acc_3_nl = ({z_out_4 , (reconstruction_error_for_l_acc_psp[1:0])})
      + ({1'b1 , (~ for_1_for_acc_6_psp_1_sva) , (~ (for_1_i_7_0_sva_4[2:0]))});
  assign reconstruction_error_for_acc_3_nl = nl_reconstruction_error_for_acc_3_nl[8:0];
  assign exit_reconstruction_error_for_sva_mx0 = MUX_s_1_2_2((~ (readslicef_9_1_8((reconstruction_error_for_acc_3_nl)))),
      (~ z_out_7_32), fsm_output[9]);
  assign nl_for_1_for_acc_6_psp_1_sva = (for_1_i_7_0_sva_4[7:3]) + 5'b1;
  assign for_1_for_acc_6_psp_1_sva = nl_for_1_for_acc_6_psp_1_sva[4:0];
  assign nl_reconstruction_error_for_l_acc_psp = ({for_1_for_acc_6_psp_1_sva , (for_1_i_7_0_sva_4[2:0])})
      + 8'b11111011;
  assign reconstruction_error_for_l_acc_psp = nl_reconstruction_error_for_l_acc_psp[7:0];
  assign nl_reconstruction_error_for_for_c_acc_psp = ({for_1_for_acc_7_psp_1_sva_1
      , (for_1_for_j_8_0_sva[2:0])}) + 9'b111111011;
  assign reconstruction_error_for_for_c_acc_psp = nl_reconstruction_error_for_for_c_acc_psp[8:0];
  assign or_tmp_30 = (fsm_output[9:6]!=4'b0000);
  assign image_net_rsci_addr_d = {z_out_1 , (for_i_7_0_sva_3[2:0])};
  assign image_net_rsci_re_d_pff = ~(((~((z_out_4[6]) | for_for_aif_oif_acc_itm_9))
      | (~(for_for_if_acc_1_tmp_5 | for_for_oif_acc_itm_8))) & (fsm_output[1]));
  assign image_floue_rsci_addr_d = {z_out_1 , (for_i_7_0_sva_3[2:0])};
  assign image_error_rsci_data_in_d = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      z_out_6, (fsm_output[2]));
  assign image_error_mux1h_nl = MUX1HOT_s_1_3_2((z_out[13]), (for_for_else_acc_itm_2[13]),
      (reconstruction_error_for_for_acc_6_sdt[13]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[7])});
  assign image_error_mux_nl = MUX_v_4_2_2((for_for_else_acc_itm_2[12:9]), (reconstruction_error_for_for_acc_6_sdt[12:9]),
      fsm_output[7]);
  assign image_error_not_2_nl = ~ (fsm_output[1]);
  assign image_error_image_error_and_nl = MUX_v_4_2_2(4'b0000, (image_error_mux_nl),
      (image_error_not_2_nl));
  assign nl_for_for_if_acc_nl = (z_out[8:0]) + conv_u2u_5_9(for_i_7_0_sva_3[7:3]);
  assign for_for_if_acc_nl = nl_for_for_if_acc_nl[8:0];
  assign image_error_mux1h_2_nl = MUX1HOT_v_9_3_2((for_for_if_acc_nl), (for_for_else_acc_itm_2[8:0]),
      (reconstruction_error_for_for_acc_6_sdt[8:0]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[7])});
  assign image_error_image_error_mux_nl = MUX_v_3_2_2((for_i_7_0_sva_3[2:0]), (reconstruction_error_for_l_sva_3[2:0]),
      fsm_output[7]);
  assign image_error_rsci_addr_d = {(image_error_mux1h_nl) , (image_error_image_error_and_nl)
      , (image_error_mux1h_2_nl) , (image_error_image_error_mux_nl)};
  assign image_error_rsci_re_d = ~ (fsm_output[7]);
  assign image_error_rsci_we_d = ~((or_11_cse & or_10_cse & (fsm_output[1])) | ((~
      for_for_if_for_for_if_and_itm_1) & (fsm_output[2])));
  assign depth_rsci_data_in_d = MUX_v_32_2_2(32'b11111111, reconstruction_error_rec_error_sva,
      z_out_7_32);
  assign depth_rsci_addr_d = {z_out_1 , (for_1_i_7_0_sva_4[2:0])};
  assign depth_rsci_we_d = ~ (fsm_output[10]);
  always @(posedge clk) begin
    if ( rst ) begin
      for_i_7_0_sva_3 <= 8'b0;
    end
    else if ( or_18_cse ) begin
      for_i_7_0_sva_3 <= MUX_v_8_2_2(8'b00000000, z_out_3, (fsm_output[4]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_j_8_0_sva_3 <= 9'b0;
      reg_return_rsc_triosy_obj_ld_cse <= 1'b0;
      for_for_else_acc_itm_2 <= 14'b0;
      for_for_if_for_for_if_and_itm_1 <= 1'b0;
      reconstruction_error_rec_error_sva <= 32'b0;
      reconstruction_error_rec_error_lpi_6 <= 32'b0;
      exit_reconstruction_error_for_for_sva_1 <= 1'b0;
      reconstruction_error_for_for_c_sva_31_9_2 <= 23'b0;
      for_1_for_slc_for_1_for_acc_7_itm_1 <= 1'b0;
      for_1_for_j_8_0_sva_4 <= 9'b0;
    end
    else begin
      for_for_j_8_0_sva_3 <= MUX_v_9_2_2(9'b000000000, for_for_j_8_0_sva_4, (not_39_nl));
      reg_return_rsc_triosy_obj_ld_cse <= (~ z_out_9_5) & (fsm_output[12]);
      for_for_else_acc_itm_2 <= nl_for_for_else_acc_itm_2[13:0];
      for_for_if_for_for_if_and_itm_1 <= or_11_cse & or_10_cse;
      reconstruction_error_rec_error_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (reconstruction_error_rec_error_mux1h_4_nl), (not_34_nl));
      reconstruction_error_rec_error_lpi_6 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (reconstruction_error_rec_error_mux1h_5_nl), (not_nl));
      exit_reconstruction_error_for_for_sva_1 <= ~ z_out_7_32;
      reconstruction_error_for_for_c_sva_31_9_2 <= MUX_v_23_2_2(23'b00000000000000000000000,
          (reconstruction_error_for_for_c_mux_nl), (not_38_nl));
      for_1_for_slc_for_1_for_acc_7_itm_1 <= z_out_2[7];
      for_1_for_j_8_0_sva_4 <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_slc_for_for_acc_7_itm <= 1'b0;
    end
    else if ( fsm_output[1] ) begin
      for_for_slc_for_for_acc_7_itm <= z_out_2[7];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_j_8_0_sva_4 <= 9'b0;
    end
    else if ( fsm_output[1] ) begin
      for_for_j_8_0_sva_4 <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_1_i_7_0_sva_4 <= 8'b0;
    end
    else if ( (fsm_output[4]) | (fsm_output[12]) ) begin
      for_1_i_7_0_sva_4 <= MUX_v_8_2_2(8'b00000000, z_out_3, (fsm_output[12]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_1_for_j_8_0_sva <= 9'b0;
    end
    else if ( (fsm_output[12]) | (fsm_output[4]) | (fsm_output[11]) ) begin
      for_1_for_j_8_0_sva <= MUX_v_9_2_2(9'b000000000, for_1_for_j_8_0_sva_4, (fsm_output[11]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_1_for_acc_6_psp_1_sva_1 <= 5'b0;
    end
    else if ( ~ or_tmp_30 ) begin
      for_1_for_acc_6_psp_1_sva_1 <= for_1_for_acc_6_psp_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reconstruction_error_for_l_sva_3 <= 32'b0;
    end
    else if ( (fsm_output[5]) | (fsm_output[9]) ) begin
      reconstruction_error_for_l_sva_3 <= MUX_v_32_2_2(({24'b0 , reconstruction_error_for_l_acc_psp}),
          z_out_8, fsm_output[9]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_1_for_acc_7_psp_1_sva_1 <= 6'b0;
    end
    else if ( ~ or_tmp_30 ) begin
      for_1_for_acc_7_psp_1_sva_1 <= nl_for_1_for_acc_7_psp_1_sva_1[5:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reconstruction_error_for_for_c_sva_8_0_2 <= 9'b0;
    end
    else if ( ~ (fsm_output[8]) ) begin
      reconstruction_error_for_for_c_sva_8_0_2 <= MUX_v_9_2_2(reconstruction_error_for_for_c_acc_psp,
          (z_out_8[8:0]), fsm_output[7]);
    end
  end
  assign not_39_nl = ~ or_18_cse;
  assign nl_for_for_else_acc_itm_2  = (z_out[13:0]) + conv_u2u_5_14(for_i_7_0_sva_3[7:3]);
  assign reconstruction_error_rec_error_mux1h_4_nl = MUX1HOT_v_32_3_2(reconstruction_error_rec_error_lpi_6,
      z_out_6, reconstruction_error_rec_error_sva, {(fsm_output[6]) , (fsm_output[8])
      , (fsm_output[9])});
  assign not_34_nl = ~ (fsm_output[5]);
  assign or_49_nl = (fsm_output[7:6]!=2'b00);
  assign reconstruction_error_rec_error_mux1h_5_nl = MUX1HOT_v_32_3_2(reconstruction_error_rec_error_lpi_6,
      z_out_6, reconstruction_error_rec_error_sva, {(or_49_nl) , (fsm_output[8])
      , (fsm_output[9])});
  assign not_nl = ~ (fsm_output[5]);
  assign reconstruction_error_for_for_c_mux_nl = MUX_v_23_2_2((z_out_8[31:9]), reconstruction_error_for_for_c_sva_31_9_2,
      fsm_output[8]);
  assign not_38_nl = ~ (fsm_output[6]);
  assign nl_for_1_for_acc_7_psp_1_sva_1  = (for_1_for_j_8_0_sva[8:3]) + 6'b1;
  assign reconstruction_error_for_for_nor_2_nl = ~((fsm_output[7]) | (fsm_output[1])
      | (fsm_output[10]));
  assign reconstruction_error_for_for_reconstruction_error_for_for_and_2_nl = MUX_v_18_2_2(18'b000000000000000000,
      (image_error_rsci_data_out_d[31:14]), (reconstruction_error_for_for_nor_2_nl));
  assign reconstruction_error_for_for_mux_3_nl = MUX_v_5_2_2((reconstruction_error_for_for_c_sva_31_9_2[4:0]),
      (image_error_rsci_data_out_d[13:9]), fsm_output[8]);
  assign reconstruction_error_for_for_nor_3_nl = ~((fsm_output[1]) | (fsm_output[10]));
  assign reconstruction_error_for_for_reconstruction_error_for_for_and_3_nl = MUX_v_5_2_2(5'b00000,
      (reconstruction_error_for_for_mux_3_nl), (reconstruction_error_for_for_nor_3_nl));
  assign reconstruction_error_for_for_mux1h_2_nl = MUX1HOT_v_9_4_2(reconstruction_error_for_for_c_sva_8_0_2,
      for_for_j_8_0_sva_3, (image_error_rsci_data_out_d[8:0]), for_1_for_j_8_0_sva,
      {(fsm_output[7]) , (fsm_output[1]) , (fsm_output[8]) , (fsm_output[10])});
  assign reconstruction_error_for_for_or_2_nl = (fsm_output[7]) | (fsm_output[1]);
  assign reconstruction_error_for_for_mux1h_3_nl = MUX1HOT_v_32_3_2(32'b11011, image_error_rsci_data_out_d,
      32'b11001, {(reconstruction_error_for_for_or_2_nl) , (fsm_output[8]) , (fsm_output[10])});
  assign nl_z_out = ({(reconstruction_error_for_for_reconstruction_error_for_for_and_2_nl)
      , (reconstruction_error_for_for_reconstruction_error_for_for_and_3_nl) , (reconstruction_error_for_for_mux1h_2_nl)})
      * (reconstruction_error_for_for_mux1h_3_nl);
  assign z_out = nl_z_out[31:0];
  assign nl_for_for_else_mul_2_nl = (for_for_j_8_0_sva_3) * 5'b11001;
  assign for_for_else_mul_2_nl = nl_for_for_else_mul_2_nl[12:0];
  assign for_for_else_mux_2_nl = MUX_v_13_2_2((for_for_else_mul_2_nl), (z_out[12:0]),
      fsm_output[10]);
  assign for_for_else_mux_3_nl = MUX_v_5_2_2((for_i_7_0_sva_3[7:3]), (for_1_i_7_0_sva_4[7:3]),
      fsm_output[10]);
  assign nl_z_out_1 = (for_for_else_mux_2_nl) + conv_u2u_5_13(for_for_else_mux_3_nl);
  assign z_out_1 = nl_z_out_1[12:0];
  assign for_for_mux1h_2_nl = MUX1HOT_v_8_3_2(8'b10110001, 8'b10110101, 8'b1111111,
      {(fsm_output[1]) , (fsm_output[10]) , (fsm_output[7])});
  assign or_60_nl = (fsm_output[1]) | (fsm_output[10]);
  assign mux_2_nl = MUX_v_7_2_2(({(~ for_1_for_acc_7_psp_1_sva_1) , (~ (for_1_for_j_8_0_sva[2]))}),
      (z_out_5[8:2]), or_60_nl);
  assign nl_z_out_2 = (for_for_mux1h_2_nl) + conv_u2u_7_8(mux_2_nl);
  assign z_out_2 = nl_z_out_2[7:0];
  assign for_mux_3_nl = MUX_v_8_2_2(for_i_7_0_sva_3, for_1_i_7_0_sva_4, fsm_output[12]);
  assign nl_z_out_3 = (for_mux_3_nl) + 8'b1;
  assign z_out_3 = nl_z_out_3[7:0];
  assign for_for_aelse_mux_4_nl = MUX_v_6_2_2((for_for_j_8_0_sva_3[8:3]), (reconstruction_error_for_l_acc_psp[7:2]),
      fsm_output[5]);
  assign nl_z_out_4 = conv_u2u_6_7(for_for_aelse_mux_4_nl) + 7'b1111111;
  assign z_out_4 = nl_z_out_4[6:0];
  assign for_for_mux_2_nl = MUX_v_9_2_2(for_for_j_8_0_sva_3, for_1_for_j_8_0_sva,
      fsm_output[10]);
  assign nl_z_out_5 = (for_for_mux_2_nl) + 9'b1;
  assign z_out_5 = nl_z_out_5[8:0];
  assign reconstruction_error_for_for_mux_4_nl = MUX_v_32_2_2(reconstruction_error_rec_error_lpi_6,
      image_floue_rsci_data_out_d, fsm_output[2]);
  assign reconstruction_error_for_for_mux_5_nl = MUX_v_32_2_2(z_out, (~ image_net_rsci_data_out_d),
      fsm_output[2]);
  assign nl_acc_5_nl = ({(reconstruction_error_for_for_mux_4_nl) , (~ (fsm_output[8]))})
      + ({(reconstruction_error_for_for_mux_5_nl) , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[32:0];
  assign z_out_6 = readslicef_33_32_1((acc_5_nl));
  assign reconstruction_error_for_reconstruction_error_for_mux_1_nl = MUX_v_32_2_2(z_out_8,
      reconstruction_error_rec_error_sva, fsm_output[10]);
  assign reconstruction_error_for_reconstruction_error_for_or_1_nl = (z_out_2[6])
      | (fsm_output[10:9]!=2'b00);
  assign nl_reconstruction_error_for_acc_8_nl = ({(~ for_1_for_acc_6_psp_1_sva_1)
      , (~ (for_1_i_7_0_sva_4[2]))}) + 6'b111111;
  assign reconstruction_error_for_acc_8_nl = nl_reconstruction_error_for_acc_8_nl[5:0];
  assign reconstruction_error_for_mux_4_nl = MUX_v_6_2_2((reconstruction_error_for_acc_8_nl),
      (z_out_2[5:0]), fsm_output[7]);
  assign reconstruction_error_for_not_13_nl = ~ (fsm_output[10]);
  assign reconstruction_error_for_reconstruction_error_for_and_1_nl = MUX_v_6_2_2(6'b000000,
      (reconstruction_error_for_mux_4_nl), (reconstruction_error_for_not_13_nl));
  assign reconstruction_error_for_mux1h_2_nl = MUX1HOT_v_2_3_2((~ (for_1_i_7_0_sva_4[1:0])),
      (~ (for_1_for_j_8_0_sva[1:0])), 2'b1, {(fsm_output[9]) , (fsm_output[7]) ,
      (fsm_output[10])});
  assign nl_reconstruction_error_for_acc_nl = conv_s2u_32_33(reconstruction_error_for_reconstruction_error_for_mux_1_nl)
      + conv_s2u_10_33({1'b1 , (reconstruction_error_for_reconstruction_error_for_or_1_nl)
      , (reconstruction_error_for_reconstruction_error_for_and_1_nl) , (reconstruction_error_for_mux1h_2_nl)});
  assign reconstruction_error_for_acc_nl = nl_reconstruction_error_for_acc_nl[32:0];
  assign z_out_7_32 = readslicef_33_1_32((reconstruction_error_for_acc_nl));
  assign reconstruction_error_for_mux_5_nl = MUX_v_32_2_2(reconstruction_error_for_l_sva_3,
      ({reconstruction_error_for_for_c_sva_31_9_2 , reconstruction_error_for_for_c_sva_8_0_2}),
      fsm_output[7]);
  assign nl_z_out_8 = (reconstruction_error_for_mux_5_nl) + 32'b1;
  assign z_out_8 = nl_z_out_8[31:0];
  assign nl_for_acc_nl = ({4'b1001 , (fsm_output[12]) , 1'b1}) + conv_u2u_5_6(z_out_3[7:3]);
  assign for_acc_nl = nl_for_acc_nl[5:0];
  assign z_out_9_5 = readslicef_6_1_5((for_acc_nl));

  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction


  function [8:0] MUX1HOT_v_9_4_2;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [3:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    MUX1HOT_v_9_4_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input [0:0] sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function [17:0] MUX_v_18_2_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [0:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_18_2_2 = result;
  end
  endfunction


  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function [7:0] readslicef_10_8_2;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_10_8_2 = tmp[7:0];
  end
  endfunction


  function [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function [31:0] readslicef_33_32_1;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_33_32_1 = tmp[31:0];
  end
  endfunction


  function [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function  [32:0] conv_s2u_10_33 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_33 = {{23{vector[9]}}, vector};
  end
  endfunction


  function  [32:0] conv_s2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_s2u_32_33 = {vector[31], vector};
  end
  endfunction


  function  [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction


  function  [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function  [8:0] conv_u2u_5_9 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_9 = {{4{1'b0}}, vector};
  end
  endfunction


  function  [12:0] conv_u2u_5_13 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_13 = {{8{1'b0}}, vector};
  end
  endfunction


  function  [13:0] conv_u2u_5_14 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_14 = {{9{1'b0}}, vector};
  end
  endfunction


  function  [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function  [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function  [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    main
// ------------------------------------------------------------------


module main (
  clk, rst, image_net_rsc_addr, image_net_rsc_re, image_net_rsc_data_out, image_net_rsc_triosy_lz,
      image_floue_rsc_addr, image_floue_rsc_re, image_floue_rsc_data_out, image_floue_rsc_triosy_lz,
      image_error_rsc_data_in, image_error_rsc_addr, image_error_rsc_re, image_error_rsc_we,
      image_error_rsc_data_out, image_error_rsc_triosy_lz, depth_rsc_data_in, depth_rsc_addr,
      depth_rsc_we, depth_rsc_triosy_lz, return_rsc_z, return_rsc_triosy_lz
);
  input clk;
  input rst;
  output [15:0] image_net_rsc_addr;
  output image_net_rsc_re;
  input [31:0] image_net_rsc_data_out;
  output image_net_rsc_triosy_lz;
  output [15:0] image_floue_rsc_addr;
  output image_floue_rsc_re;
  input [31:0] image_floue_rsc_data_out;
  output image_floue_rsc_triosy_lz;
  output [31:0] image_error_rsc_data_in;
  output [16:0] image_error_rsc_addr;
  output image_error_rsc_re;
  output image_error_rsc_we;
  input [31:0] image_error_rsc_data_out;
  output image_error_rsc_triosy_lz;
  output [31:0] depth_rsc_data_in;
  output [15:0] depth_rsc_addr;
  output depth_rsc_we;
  output depth_rsc_triosy_lz;
  output [31:0] return_rsc_z;
  output return_rsc_triosy_lz;


  // Interconnect Declarations
  wire [15:0] image_net_rsci_addr_d;
  wire [31:0] image_net_rsci_data_out_d;
  wire [15:0] image_floue_rsci_addr_d;
  wire [31:0] image_floue_rsci_data_out_d;
  wire [31:0] image_error_rsci_data_in_d;
  wire [16:0] image_error_rsci_addr_d;
  wire image_error_rsci_re_d;
  wire image_error_rsci_we_d;
  wire [31:0] image_error_rsci_data_out_d;
  wire [31:0] depth_rsci_data_in_d;
  wire [15:0] depth_rsci_addr_d;
  wire depth_rsci_we_d;
  wire image_net_rsci_re_d_iff;


  // Interconnect Declarations for Component Instantiations 
  ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rport_3_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
      image_net_rsci (
      .data_out(image_net_rsc_data_out),
      .re(image_net_rsc_re),
      .addr(image_net_rsc_addr),
      .addr_d(image_net_rsci_addr_d),
      .re_d(image_net_rsci_re_d_iff),
      .data_out_d(image_net_rsci_data_out_d)
    );
  ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rport_4_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
      image_floue_rsci (
      .data_out(image_floue_rsc_data_out),
      .re(image_floue_rsc_re),
      .addr(image_floue_rsc_addr),
      .addr_d(image_floue_rsci_addr_d),
      .re_d(image_net_rsci_re_d_iff),
      .data_out_d(image_floue_rsci_data_out_d)
    );
  ram_Xilinx_KINTEX_7_3_RAMSB_singleport_rwport_5_68256_32_17_0_1_0_0_0_1_1_1_0_68256_32_1_gen
      image_error_rsci (
      .data_out(image_error_rsc_data_out),
      .we(image_error_rsc_we),
      .re(image_error_rsc_re),
      .addr(image_error_rsc_addr),
      .data_in(image_error_rsc_data_in),
      .data_in_d(image_error_rsci_data_in_d),
      .addr_d(image_error_rsci_addr_d),
      .re_d(image_error_rsci_re_d),
      .we_d(image_error_rsci_we_d),
      .data_out_d(image_error_rsci_data_out_d)
    );
  ram_Xilinx_KINTEX_7_3_RAMSB_singleport_wport_6_60000_32_16_0_1_0_0_0_1_1_1_0_60000_32_1_gen
      depth_rsci (
      .we(depth_rsc_we),
      .addr(depth_rsc_addr),
      .data_in(depth_rsc_data_in),
      .data_in_d(depth_rsci_data_in_d),
      .addr_d(depth_rsci_addr_d),
      .we_d(depth_rsci_we_d)
    );
  main_core main_core_inst (
      .clk(clk),
      .rst(rst),
      .image_net_rsc_triosy_lz(image_net_rsc_triosy_lz),
      .image_floue_rsc_triosy_lz(image_floue_rsc_triosy_lz),
      .image_error_rsc_triosy_lz(image_error_rsc_triosy_lz),
      .depth_rsc_triosy_lz(depth_rsc_triosy_lz),
      .return_rsc_z(return_rsc_z),
      .return_rsc_triosy_lz(return_rsc_triosy_lz),
      .image_net_rsci_addr_d(image_net_rsci_addr_d),
      .image_net_rsci_data_out_d(image_net_rsci_data_out_d),
      .image_floue_rsci_addr_d(image_floue_rsci_addr_d),
      .image_floue_rsci_data_out_d(image_floue_rsci_data_out_d),
      .image_error_rsci_data_in_d(image_error_rsci_data_in_d),
      .image_error_rsci_addr_d(image_error_rsci_addr_d),
      .image_error_rsci_re_d(image_error_rsci_re_d),
      .image_error_rsci_we_d(image_error_rsci_we_d),
      .image_error_rsci_data_out_d(image_error_rsci_data_out_d),
      .depth_rsci_data_in_d(depth_rsci_data_in_d),
      .depth_rsci_addr_d(depth_rsci_addr_d),
      .depth_rsci_we_d(depth_rsci_we_d),
      .image_net_rsci_re_d_pff(image_net_rsci_re_d_iff)
    );
endmodule



