//
// Verilog description for cell main, 
// Tue Jan 16 15:04:54 2018
//
// Precision RTL Synthesis, 2014a.1_64-bit//


module main ( clk, rst, image_net_rsc_addr, image_net_rsc_re, 
              image_net_rsc_data_out, image_net_rsc_triosy_lz, 
              image_floue_rsc_addr, image_floue_rsc_re, image_floue_rsc_data_out, 
              image_floue_rsc_triosy_lz, image_error_rsc_data_in, 
              image_error_rsc_addr, image_error_rsc_re, image_error_rsc_we, 
              image_error_rsc_data_out, image_error_rsc_triosy_lz, 
              depth_rsc_data_in, depth_rsc_addr, depth_rsc_we, 
              depth_rsc_triosy_lz, return_rsc_z, return_rsc_triosy_lz ) ;

    input clk ;
    input rst ;
    output [15:0]image_net_rsc_addr ;
    output image_net_rsc_re ;
    input [31:0]image_net_rsc_data_out ;
    output image_net_rsc_triosy_lz ;
    output [15:0]image_floue_rsc_addr ;
    output image_floue_rsc_re ;
    input [31:0]image_floue_rsc_data_out ;
    output image_floue_rsc_triosy_lz ;
    output [31:0]image_error_rsc_data_in ;
    output [16:0]image_error_rsc_addr ;
    output image_error_rsc_re ;
    output image_error_rsc_we ;
    input [31:0]image_error_rsc_data_out ;
    output image_error_rsc_triosy_lz ;
    output [31:0]depth_rsc_data_in ;
    output [15:0]depth_rsc_addr ;
    output depth_rsc_we ;
    output depth_rsc_triosy_lz ;
    output [31:0]return_rsc_z ;
    output return_rsc_triosy_lz ;

    wire [15:0]image_net_rsc_addr_1_0;
    wire image_net_rsc_triosy_lz_1_0;
    wire [2:0]depth_rsc_addr_1_0;
    wire clk_int;
    wire rst_int;
    wire [31:0]image_net_rsc_data_out_int;
    wire [31:0]image_floue_rsc_data_out_int;
    wire [31:0]image_error_rsc_data_out_int;
    wire \main_core_inst_fsm_output(10)  ;
    wire \main_core_inst_z_out(8)  , \main_core_inst_z_out(7)  , 
         \main_core_inst_z_out(6)  , \main_core_inst_z_out(5)  , 
         \main_core_inst_z_out(4)  , \main_core_inst_z_out(3)  , 
         \main_core_inst_z_out(2)  , \main_core_inst_z_out(1)  , 
         \main_core_inst_z_out(0)  ;
    wire \main_core_inst_for_for_mux1h_2_nl(1)  ;
    wire image_error_rsc_re_1_0, depth_rsc_we_1_0, nx18058z10, nx18058z1, 
         nx18058z2, nx18058z3, nx18058z4, nx18058z5, nx18058z6, nx18058z7, 
         nx18058z8, nx18058z9, nx7721z1, nx56118z1, nx55121z1, nx53125z1, 
         nx52128z1, nx51131z1, nx50134z1, nx49137z1, nx48140z1, nx47143z1, 
         nx46146z1, nx45149z1, nx44152z1, nx42156z1, nx41159z1, nx40162z1, 
         nx39165z1, nx38168z1, nx37171z1, nx36174z1, nx35177z1, nx34180z1, 
         nx33183z1, nx28511z1, nx27514z1, nx26517z1, nx25520z1, nx24523z1, 
         nx23526z1, nx22529z1, nx21532z1, nx20535z1, nx19538z1, nx16900z1, 
         nx17897z1, nx18894z1, nx19891z1, nx20888z1, nx21885z1, nx22882z1, 
         nx53646z1, nx54643z1, nx55640z1, nx56637z1, nx57634z1, nx58631z1, 
         nx59628z1, nx60625z1, nx61622z1, nx62619z1, nx51351z1, nx32759z1, 
         nx31762z1, nx29766z1, nx28769z1, nx27772z1, nx26775z1, nx25778z1, 
         nx24781z1, nx23784z1, nx22787z1, nx21790z1, nx20793z1, nx18797z1, 
         nx17800z1, nx16803z1, nx15806z1, nx14809z1, nx13812z1, nx12815z1, 
         nx11818z1, nx10821z1, nx9824z1, nx51444z1, nx52441z1, nx53438z1, 
         nx54435z1, nx55432z1, nx56429z1, nx57426z1, nx58423z1, nx59420z1, 
         nx60417z1, nx18058z11;



    OBUF return_rsc_triosy_lz_obuf (.O (return_rsc_triosy_lz), .I (
         image_net_rsc_triosy_lz_1_0)) ;
    OBUF \return_rsc_z_obuf(0)  (.O (return_rsc_z[0]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(1)  (.O (return_rsc_z[1]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(2)  (.O (return_rsc_z[2]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(3)  (.O (return_rsc_z[3]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(4)  (.O (return_rsc_z[4]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(5)  (.O (return_rsc_z[5]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(6)  (.O (return_rsc_z[6]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(7)  (.O (return_rsc_z[7]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(8)  (.O (return_rsc_z[8]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(9)  (.O (return_rsc_z[9]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(10)  (.O (return_rsc_z[10]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(11)  (.O (return_rsc_z[11]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(12)  (.O (return_rsc_z[12]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(13)  (.O (return_rsc_z[13]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(14)  (.O (return_rsc_z[14]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(15)  (.O (return_rsc_z[15]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(16)  (.O (return_rsc_z[16]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(17)  (.O (return_rsc_z[17]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(18)  (.O (return_rsc_z[18]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(19)  (.O (return_rsc_z[19]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(20)  (.O (return_rsc_z[20]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(21)  (.O (return_rsc_z[21]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(22)  (.O (return_rsc_z[22]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(23)  (.O (return_rsc_z[23]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(24)  (.O (return_rsc_z[24]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(25)  (.O (return_rsc_z[25]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(26)  (.O (return_rsc_z[26]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(27)  (.O (return_rsc_z[27]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(28)  (.O (return_rsc_z[28]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(29)  (.O (return_rsc_z[29]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(30)  (.O (return_rsc_z[30]), .I (nx18058z10)) ;
    OBUF \return_rsc_z_obuf(31)  (.O (return_rsc_z[31]), .I (nx18058z10)) ;
    OBUF depth_rsc_triosy_lz_obuf (.O (depth_rsc_triosy_lz), .I (
         image_net_rsc_triosy_lz_1_0)) ;
    OBUF depth_rsc_we_obuf (.O (depth_rsc_we), .I (depth_rsc_we_1_0)) ;
    OBUF \depth_rsc_addr_obuf(0)  (.O (depth_rsc_addr[0]), .I (
         depth_rsc_addr_1_0[0])) ;
    OBUF \depth_rsc_addr_obuf(1)  (.O (depth_rsc_addr[1]), .I (
         depth_rsc_addr_1_0[1])) ;
    OBUF \depth_rsc_addr_obuf(2)  (.O (depth_rsc_addr[2]), .I (
         depth_rsc_addr_1_0[2])) ;
    OBUF \depth_rsc_addr_obuf(3)  (.O (depth_rsc_addr[3]), .I (
         image_net_rsc_addr_1_0[3])) ;
    OBUF \depth_rsc_addr_obuf(4)  (.O (depth_rsc_addr[4]), .I (
         image_net_rsc_addr_1_0[4])) ;
    OBUF \depth_rsc_addr_obuf(5)  (.O (depth_rsc_addr[5]), .I (
         image_net_rsc_addr_1_0[5])) ;
    OBUF \depth_rsc_addr_obuf(6)  (.O (depth_rsc_addr[6]), .I (
         image_net_rsc_addr_1_0[6])) ;
    OBUF \depth_rsc_addr_obuf(7)  (.O (depth_rsc_addr[7]), .I (
         image_net_rsc_addr_1_0[7])) ;
    OBUF \depth_rsc_addr_obuf(8)  (.O (depth_rsc_addr[8]), .I (
         image_net_rsc_addr_1_0[8])) ;
    OBUF \depth_rsc_addr_obuf(9)  (.O (depth_rsc_addr[9]), .I (
         image_net_rsc_addr_1_0[9])) ;
    OBUF \depth_rsc_addr_obuf(10)  (.O (depth_rsc_addr[10]), .I (
         image_net_rsc_addr_1_0[10])) ;
    OBUF \depth_rsc_addr_obuf(11)  (.O (depth_rsc_addr[11]), .I (
         image_net_rsc_addr_1_0[11])) ;
    OBUF \depth_rsc_addr_obuf(12)  (.O (depth_rsc_addr[12]), .I (
         image_net_rsc_addr_1_0[12])) ;
    OBUF \depth_rsc_addr_obuf(13)  (.O (depth_rsc_addr[13]), .I (
         image_net_rsc_addr_1_0[13])) ;
    OBUF \depth_rsc_addr_obuf(14)  (.O (depth_rsc_addr[14]), .I (
         image_net_rsc_addr_1_0[14])) ;
    OBUF \depth_rsc_addr_obuf(15)  (.O (depth_rsc_addr[15]), .I (
         image_net_rsc_addr_1_0[15])) ;
    OBUF \depth_rsc_data_in_obuf(0)  (.O (depth_rsc_data_in[0]), .I (nx60417z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(1)  (.O (depth_rsc_data_in[1]), .I (nx59420z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(2)  (.O (depth_rsc_data_in[2]), .I (nx58423z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(3)  (.O (depth_rsc_data_in[3]), .I (nx57426z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(4)  (.O (depth_rsc_data_in[4]), .I (nx56429z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(5)  (.O (depth_rsc_data_in[5]), .I (nx55432z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(6)  (.O (depth_rsc_data_in[6]), .I (nx54435z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(7)  (.O (depth_rsc_data_in[7]), .I (nx53438z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(8)  (.O (depth_rsc_data_in[8]), .I (nx52441z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(9)  (.O (depth_rsc_data_in[9]), .I (nx51444z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(10)  (.O (depth_rsc_data_in[10]), .I (nx9824z1)
         ) ;
    OBUF \depth_rsc_data_in_obuf(11)  (.O (depth_rsc_data_in[11]), .I (nx10821z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(12)  (.O (depth_rsc_data_in[12]), .I (nx11818z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(13)  (.O (depth_rsc_data_in[13]), .I (nx12815z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(14)  (.O (depth_rsc_data_in[14]), .I (nx13812z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(15)  (.O (depth_rsc_data_in[15]), .I (nx14809z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(16)  (.O (depth_rsc_data_in[16]), .I (nx15806z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(17)  (.O (depth_rsc_data_in[17]), .I (nx16803z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(18)  (.O (depth_rsc_data_in[18]), .I (nx17800z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(19)  (.O (depth_rsc_data_in[19]), .I (nx18797z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(20)  (.O (depth_rsc_data_in[20]), .I (nx20793z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(21)  (.O (depth_rsc_data_in[21]), .I (nx21790z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(22)  (.O (depth_rsc_data_in[22]), .I (nx22787z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(23)  (.O (depth_rsc_data_in[23]), .I (nx23784z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(24)  (.O (depth_rsc_data_in[24]), .I (nx24781z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(25)  (.O (depth_rsc_data_in[25]), .I (nx25778z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(26)  (.O (depth_rsc_data_in[26]), .I (nx26775z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(27)  (.O (depth_rsc_data_in[27]), .I (nx27772z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(28)  (.O (depth_rsc_data_in[28]), .I (nx28769z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(29)  (.O (depth_rsc_data_in[29]), .I (nx29766z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(30)  (.O (depth_rsc_data_in[30]), .I (nx31762z1
         )) ;
    OBUF \depth_rsc_data_in_obuf(31)  (.O (depth_rsc_data_in[31]), .I (nx32759z1
         )) ;
    OBUF image_error_rsc_triosy_lz_obuf (.O (image_error_rsc_triosy_lz), .I (
         image_net_rsc_triosy_lz_1_0)) ;
    OBUF image_error_rsc_we_obuf (.O (image_error_rsc_we), .I (nx51351z1)) ;
    OBUF image_error_rsc_re_obuf (.O (image_error_rsc_re), .I (
         image_error_rsc_re_1_0)) ;
    OBUF \image_error_rsc_addr_obuf(0)  (.O (image_error_rsc_addr[0]), .I (
         nx62619z1)) ;
    OBUF \image_error_rsc_addr_obuf(1)  (.O (image_error_rsc_addr[1]), .I (
         nx61622z1)) ;
    OBUF \image_error_rsc_addr_obuf(2)  (.O (image_error_rsc_addr[2]), .I (
         nx60625z1)) ;
    OBUF \image_error_rsc_addr_obuf(3)  (.O (image_error_rsc_addr[3]), .I (
         nx59628z1)) ;
    OBUF \image_error_rsc_addr_obuf(4)  (.O (image_error_rsc_addr[4]), .I (
         nx58631z1)) ;
    OBUF \image_error_rsc_addr_obuf(5)  (.O (image_error_rsc_addr[5]), .I (
         nx57634z1)) ;
    OBUF \image_error_rsc_addr_obuf(6)  (.O (image_error_rsc_addr[6]), .I (
         nx56637z1)) ;
    OBUF \image_error_rsc_addr_obuf(7)  (.O (image_error_rsc_addr[7]), .I (
         nx55640z1)) ;
    OBUF \image_error_rsc_addr_obuf(8)  (.O (image_error_rsc_addr[8]), .I (
         nx54643z1)) ;
    OBUF \image_error_rsc_addr_obuf(9)  (.O (image_error_rsc_addr[9]), .I (
         nx53646z1)) ;
    OBUF \image_error_rsc_addr_obuf(10)  (.O (image_error_rsc_addr[10]), .I (
         nx22882z1)) ;
    OBUF \image_error_rsc_addr_obuf(11)  (.O (image_error_rsc_addr[11]), .I (
         nx21885z1)) ;
    OBUF \image_error_rsc_addr_obuf(12)  (.O (image_error_rsc_addr[12]), .I (
         nx20888z1)) ;
    OBUF \image_error_rsc_addr_obuf(13)  (.O (image_error_rsc_addr[13]), .I (
         nx19891z1)) ;
    OBUF \image_error_rsc_addr_obuf(14)  (.O (image_error_rsc_addr[14]), .I (
         nx18894z1)) ;
    OBUF \image_error_rsc_addr_obuf(15)  (.O (image_error_rsc_addr[15]), .I (
         nx17897z1)) ;
    OBUF \image_error_rsc_addr_obuf(16)  (.O (image_error_rsc_addr[16]), .I (
         nx16900z1)) ;
    OBUF \image_error_rsc_data_in_obuf(0)  (.O (image_error_rsc_data_in[0]), .I (
         nx19538z1)) ;
    OBUF \image_error_rsc_data_in_obuf(1)  (.O (image_error_rsc_data_in[1]), .I (
         nx20535z1)) ;
    OBUF \image_error_rsc_data_in_obuf(2)  (.O (image_error_rsc_data_in[2]), .I (
         nx21532z1)) ;
    OBUF \image_error_rsc_data_in_obuf(3)  (.O (image_error_rsc_data_in[3]), .I (
         nx22529z1)) ;
    OBUF \image_error_rsc_data_in_obuf(4)  (.O (image_error_rsc_data_in[4]), .I (
         nx23526z1)) ;
    OBUF \image_error_rsc_data_in_obuf(5)  (.O (image_error_rsc_data_in[5]), .I (
         nx24523z1)) ;
    OBUF \image_error_rsc_data_in_obuf(6)  (.O (image_error_rsc_data_in[6]), .I (
         nx25520z1)) ;
    OBUF \image_error_rsc_data_in_obuf(7)  (.O (image_error_rsc_data_in[7]), .I (
         nx26517z1)) ;
    OBUF \image_error_rsc_data_in_obuf(8)  (.O (image_error_rsc_data_in[8]), .I (
         nx27514z1)) ;
    OBUF \image_error_rsc_data_in_obuf(9)  (.O (image_error_rsc_data_in[9]), .I (
         nx28511z1)) ;
    OBUF \image_error_rsc_data_in_obuf(10)  (.O (image_error_rsc_data_in[10]), .I (
         nx33183z1)) ;
    OBUF \image_error_rsc_data_in_obuf(11)  (.O (image_error_rsc_data_in[11]), .I (
         nx34180z1)) ;
    OBUF \image_error_rsc_data_in_obuf(12)  (.O (image_error_rsc_data_in[12]), .I (
         nx35177z1)) ;
    OBUF \image_error_rsc_data_in_obuf(13)  (.O (image_error_rsc_data_in[13]), .I (
         nx36174z1)) ;
    OBUF \image_error_rsc_data_in_obuf(14)  (.O (image_error_rsc_data_in[14]), .I (
         nx37171z1)) ;
    OBUF \image_error_rsc_data_in_obuf(15)  (.O (image_error_rsc_data_in[15]), .I (
         nx38168z1)) ;
    OBUF \image_error_rsc_data_in_obuf(16)  (.O (image_error_rsc_data_in[16]), .I (
         nx39165z1)) ;
    OBUF \image_error_rsc_data_in_obuf(17)  (.O (image_error_rsc_data_in[17]), .I (
         nx40162z1)) ;
    OBUF \image_error_rsc_data_in_obuf(18)  (.O (image_error_rsc_data_in[18]), .I (
         nx41159z1)) ;
    OBUF \image_error_rsc_data_in_obuf(19)  (.O (image_error_rsc_data_in[19]), .I (
         nx42156z1)) ;
    OBUF \image_error_rsc_data_in_obuf(20)  (.O (image_error_rsc_data_in[20]), .I (
         nx44152z1)) ;
    OBUF \image_error_rsc_data_in_obuf(21)  (.O (image_error_rsc_data_in[21]), .I (
         nx45149z1)) ;
    OBUF \image_error_rsc_data_in_obuf(22)  (.O (image_error_rsc_data_in[22]), .I (
         nx46146z1)) ;
    OBUF \image_error_rsc_data_in_obuf(23)  (.O (image_error_rsc_data_in[23]), .I (
         nx47143z1)) ;
    OBUF \image_error_rsc_data_in_obuf(24)  (.O (image_error_rsc_data_in[24]), .I (
         nx48140z1)) ;
    OBUF \image_error_rsc_data_in_obuf(25)  (.O (image_error_rsc_data_in[25]), .I (
         nx49137z1)) ;
    OBUF \image_error_rsc_data_in_obuf(26)  (.O (image_error_rsc_data_in[26]), .I (
         nx50134z1)) ;
    OBUF \image_error_rsc_data_in_obuf(27)  (.O (image_error_rsc_data_in[27]), .I (
         nx51131z1)) ;
    OBUF \image_error_rsc_data_in_obuf(28)  (.O (image_error_rsc_data_in[28]), .I (
         nx52128z1)) ;
    OBUF \image_error_rsc_data_in_obuf(29)  (.O (image_error_rsc_data_in[29]), .I (
         nx53125z1)) ;
    OBUF \image_error_rsc_data_in_obuf(30)  (.O (image_error_rsc_data_in[30]), .I (
         nx55121z1)) ;
    OBUF \image_error_rsc_data_in_obuf(31)  (.O (image_error_rsc_data_in[31]), .I (
         nx56118z1)) ;
    OBUF image_floue_rsc_triosy_lz_obuf (.O (image_floue_rsc_triosy_lz), .I (
         image_net_rsc_triosy_lz_1_0)) ;
    OBUF image_floue_rsc_re_obuf (.O (image_floue_rsc_re), .I (nx7721z1)) ;
    OBUF \image_floue_rsc_addr_obuf(0)  (.O (image_floue_rsc_addr[0]), .I (
         image_net_rsc_addr_1_0[0])) ;
    OBUF \image_floue_rsc_addr_obuf(1)  (.O (image_floue_rsc_addr[1]), .I (
         image_net_rsc_addr_1_0[1])) ;
    OBUF \image_floue_rsc_addr_obuf(2)  (.O (image_floue_rsc_addr[2]), .I (
         image_net_rsc_addr_1_0[2])) ;
    OBUF \image_floue_rsc_addr_obuf(3)  (.O (image_floue_rsc_addr[3]), .I (
         image_net_rsc_addr_1_0[3])) ;
    OBUF \image_floue_rsc_addr_obuf(4)  (.O (image_floue_rsc_addr[4]), .I (
         image_net_rsc_addr_1_0[4])) ;
    OBUF \image_floue_rsc_addr_obuf(5)  (.O (image_floue_rsc_addr[5]), .I (
         image_net_rsc_addr_1_0[5])) ;
    OBUF \image_floue_rsc_addr_obuf(6)  (.O (image_floue_rsc_addr[6]), .I (
         image_net_rsc_addr_1_0[6])) ;
    OBUF \image_floue_rsc_addr_obuf(7)  (.O (image_floue_rsc_addr[7]), .I (
         image_net_rsc_addr_1_0[7])) ;
    OBUF \image_floue_rsc_addr_obuf(8)  (.O (image_floue_rsc_addr[8]), .I (
         image_net_rsc_addr_1_0[8])) ;
    OBUF \image_floue_rsc_addr_obuf(9)  (.O (image_floue_rsc_addr[9]), .I (
         image_net_rsc_addr_1_0[9])) ;
    OBUF \image_floue_rsc_addr_obuf(10)  (.O (image_floue_rsc_addr[10]), .I (
         image_net_rsc_addr_1_0[10])) ;
    OBUF \image_floue_rsc_addr_obuf(11)  (.O (image_floue_rsc_addr[11]), .I (
         image_net_rsc_addr_1_0[11])) ;
    OBUF \image_floue_rsc_addr_obuf(12)  (.O (image_floue_rsc_addr[12]), .I (
         image_net_rsc_addr_1_0[12])) ;
    OBUF \image_floue_rsc_addr_obuf(13)  (.O (image_floue_rsc_addr[13]), .I (
         image_net_rsc_addr_1_0[13])) ;
    OBUF \image_floue_rsc_addr_obuf(14)  (.O (image_floue_rsc_addr[14]), .I (
         image_net_rsc_addr_1_0[14])) ;
    OBUF \image_floue_rsc_addr_obuf(15)  (.O (image_floue_rsc_addr[15]), .I (
         image_net_rsc_addr_1_0[15])) ;
    OBUF image_net_rsc_triosy_lz_obuf (.O (image_net_rsc_triosy_lz), .I (
         image_net_rsc_triosy_lz_1_0)) ;
    OBUF image_net_rsc_re_obuf (.O (image_net_rsc_re), .I (nx7721z1)) ;
    OBUF \image_net_rsc_addr_obuf(0)  (.O (image_net_rsc_addr[0]), .I (
         image_net_rsc_addr_1_0[0])) ;
    OBUF \image_net_rsc_addr_obuf(1)  (.O (image_net_rsc_addr[1]), .I (
         image_net_rsc_addr_1_0[1])) ;
    OBUF \image_net_rsc_addr_obuf(2)  (.O (image_net_rsc_addr[2]), .I (
         image_net_rsc_addr_1_0[2])) ;
    OBUF \image_net_rsc_addr_obuf(3)  (.O (image_net_rsc_addr[3]), .I (
         image_net_rsc_addr_1_0[3])) ;
    OBUF \image_net_rsc_addr_obuf(4)  (.O (image_net_rsc_addr[4]), .I (
         image_net_rsc_addr_1_0[4])) ;
    OBUF \image_net_rsc_addr_obuf(5)  (.O (image_net_rsc_addr[5]), .I (
         image_net_rsc_addr_1_0[5])) ;
    OBUF \image_net_rsc_addr_obuf(6)  (.O (image_net_rsc_addr[6]), .I (
         image_net_rsc_addr_1_0[6])) ;
    OBUF \image_net_rsc_addr_obuf(7)  (.O (image_net_rsc_addr[7]), .I (
         image_net_rsc_addr_1_0[7])) ;
    OBUF \image_net_rsc_addr_obuf(8)  (.O (image_net_rsc_addr[8]), .I (
         image_net_rsc_addr_1_0[8])) ;
    OBUF \image_net_rsc_addr_obuf(9)  (.O (image_net_rsc_addr[9]), .I (
         image_net_rsc_addr_1_0[9])) ;
    OBUF \image_net_rsc_addr_obuf(10)  (.O (image_net_rsc_addr[10]), .I (
         image_net_rsc_addr_1_0[10])) ;
    OBUF \image_net_rsc_addr_obuf(11)  (.O (image_net_rsc_addr[11]), .I (
         image_net_rsc_addr_1_0[11])) ;
    OBUF \image_net_rsc_addr_obuf(12)  (.O (image_net_rsc_addr[12]), .I (
         image_net_rsc_addr_1_0[12])) ;
    OBUF \image_net_rsc_addr_obuf(13)  (.O (image_net_rsc_addr[13]), .I (
         image_net_rsc_addr_1_0[13])) ;
    OBUF \image_net_rsc_addr_obuf(14)  (.O (image_net_rsc_addr[14]), .I (
         image_net_rsc_addr_1_0[14])) ;
    OBUF \image_net_rsc_addr_obuf(15)  (.O (image_net_rsc_addr[15]), .I (
         image_net_rsc_addr_1_0[15])) ;
    IBUF \image_error_rsc_data_out_ibuf(0)  (.O (image_error_rsc_data_out_int[0]
         ), .I (image_error_rsc_data_out[0])) ;
    IBUF \image_error_rsc_data_out_ibuf(1)  (.O (image_error_rsc_data_out_int[1]
         ), .I (image_error_rsc_data_out[1])) ;
    IBUF \image_error_rsc_data_out_ibuf(2)  (.O (image_error_rsc_data_out_int[2]
         ), .I (image_error_rsc_data_out[2])) ;
    IBUF \image_error_rsc_data_out_ibuf(3)  (.O (image_error_rsc_data_out_int[3]
         ), .I (image_error_rsc_data_out[3])) ;
    IBUF \image_error_rsc_data_out_ibuf(4)  (.O (image_error_rsc_data_out_int[4]
         ), .I (image_error_rsc_data_out[4])) ;
    IBUF \image_error_rsc_data_out_ibuf(5)  (.O (image_error_rsc_data_out_int[5]
         ), .I (image_error_rsc_data_out[5])) ;
    IBUF \image_error_rsc_data_out_ibuf(6)  (.O (image_error_rsc_data_out_int[6]
         ), .I (image_error_rsc_data_out[6])) ;
    IBUF \image_error_rsc_data_out_ibuf(7)  (.O (image_error_rsc_data_out_int[7]
         ), .I (image_error_rsc_data_out[7])) ;
    IBUF \image_error_rsc_data_out_ibuf(8)  (.O (image_error_rsc_data_out_int[8]
         ), .I (image_error_rsc_data_out[8])) ;
    IBUF \image_error_rsc_data_out_ibuf(9)  (.O (image_error_rsc_data_out_int[9]
         ), .I (image_error_rsc_data_out[9])) ;
    IBUF \image_error_rsc_data_out_ibuf(10)  (.O (
         image_error_rsc_data_out_int[10]), .I (image_error_rsc_data_out[10])) ;
    IBUF \image_error_rsc_data_out_ibuf(11)  (.O (
         image_error_rsc_data_out_int[11]), .I (image_error_rsc_data_out[11])) ;
    IBUF \image_error_rsc_data_out_ibuf(12)  (.O (
         image_error_rsc_data_out_int[12]), .I (image_error_rsc_data_out[12])) ;
    IBUF \image_error_rsc_data_out_ibuf(13)  (.O (
         image_error_rsc_data_out_int[13]), .I (image_error_rsc_data_out[13])) ;
    IBUF \image_error_rsc_data_out_ibuf(14)  (.O (
         image_error_rsc_data_out_int[14]), .I (image_error_rsc_data_out[14])) ;
    IBUF \image_error_rsc_data_out_ibuf(15)  (.O (
         image_error_rsc_data_out_int[15]), .I (image_error_rsc_data_out[15])) ;
    IBUF \image_error_rsc_data_out_ibuf(16)  (.O (
         image_error_rsc_data_out_int[16]), .I (image_error_rsc_data_out[16])) ;
    IBUF \image_error_rsc_data_out_ibuf(17)  (.O (
         image_error_rsc_data_out_int[17]), .I (image_error_rsc_data_out[17])) ;
    IBUF \image_error_rsc_data_out_ibuf(18)  (.O (
         image_error_rsc_data_out_int[18]), .I (image_error_rsc_data_out[18])) ;
    IBUF \image_error_rsc_data_out_ibuf(19)  (.O (
         image_error_rsc_data_out_int[19]), .I (image_error_rsc_data_out[19])) ;
    IBUF \image_error_rsc_data_out_ibuf(20)  (.O (
         image_error_rsc_data_out_int[20]), .I (image_error_rsc_data_out[20])) ;
    IBUF \image_error_rsc_data_out_ibuf(21)  (.O (
         image_error_rsc_data_out_int[21]), .I (image_error_rsc_data_out[21])) ;
    IBUF \image_error_rsc_data_out_ibuf(22)  (.O (
         image_error_rsc_data_out_int[22]), .I (image_error_rsc_data_out[22])) ;
    IBUF \image_error_rsc_data_out_ibuf(23)  (.O (
         image_error_rsc_data_out_int[23]), .I (image_error_rsc_data_out[23])) ;
    IBUF \image_error_rsc_data_out_ibuf(24)  (.O (
         image_error_rsc_data_out_int[24]), .I (image_error_rsc_data_out[24])) ;
    IBUF \image_error_rsc_data_out_ibuf(25)  (.O (
         image_error_rsc_data_out_int[25]), .I (image_error_rsc_data_out[25])) ;
    IBUF \image_error_rsc_data_out_ibuf(26)  (.O (
         image_error_rsc_data_out_int[26]), .I (image_error_rsc_data_out[26])) ;
    IBUF \image_error_rsc_data_out_ibuf(27)  (.O (
         image_error_rsc_data_out_int[27]), .I (image_error_rsc_data_out[27])) ;
    IBUF \image_error_rsc_data_out_ibuf(28)  (.O (
         image_error_rsc_data_out_int[28]), .I (image_error_rsc_data_out[28])) ;
    IBUF \image_error_rsc_data_out_ibuf(29)  (.O (
         image_error_rsc_data_out_int[29]), .I (image_error_rsc_data_out[29])) ;
    IBUF \image_error_rsc_data_out_ibuf(30)  (.O (
         image_error_rsc_data_out_int[30]), .I (image_error_rsc_data_out[30])) ;
    IBUF \image_error_rsc_data_out_ibuf(31)  (.O (
         image_error_rsc_data_out_int[31]), .I (image_error_rsc_data_out[31])) ;
    IBUF \image_floue_rsc_data_out_ibuf(0)  (.O (image_floue_rsc_data_out_int[0]
         ), .I (image_floue_rsc_data_out[0])) ;
    IBUF \image_floue_rsc_data_out_ibuf(1)  (.O (image_floue_rsc_data_out_int[1]
         ), .I (image_floue_rsc_data_out[1])) ;
    IBUF \image_floue_rsc_data_out_ibuf(2)  (.O (image_floue_rsc_data_out_int[2]
         ), .I (image_floue_rsc_data_out[2])) ;
    IBUF \image_floue_rsc_data_out_ibuf(3)  (.O (image_floue_rsc_data_out_int[3]
         ), .I (image_floue_rsc_data_out[3])) ;
    IBUF \image_floue_rsc_data_out_ibuf(4)  (.O (image_floue_rsc_data_out_int[4]
         ), .I (image_floue_rsc_data_out[4])) ;
    IBUF \image_floue_rsc_data_out_ibuf(5)  (.O (image_floue_rsc_data_out_int[5]
         ), .I (image_floue_rsc_data_out[5])) ;
    IBUF \image_floue_rsc_data_out_ibuf(6)  (.O (image_floue_rsc_data_out_int[6]
         ), .I (image_floue_rsc_data_out[6])) ;
    IBUF \image_floue_rsc_data_out_ibuf(7)  (.O (image_floue_rsc_data_out_int[7]
         ), .I (image_floue_rsc_data_out[7])) ;
    IBUF \image_floue_rsc_data_out_ibuf(8)  (.O (image_floue_rsc_data_out_int[8]
         ), .I (image_floue_rsc_data_out[8])) ;
    IBUF \image_floue_rsc_data_out_ibuf(9)  (.O (image_floue_rsc_data_out_int[9]
         ), .I (image_floue_rsc_data_out[9])) ;
    IBUF \image_floue_rsc_data_out_ibuf(10)  (.O (
         image_floue_rsc_data_out_int[10]), .I (image_floue_rsc_data_out[10])) ;
    IBUF \image_floue_rsc_data_out_ibuf(11)  (.O (
         image_floue_rsc_data_out_int[11]), .I (image_floue_rsc_data_out[11])) ;
    IBUF \image_floue_rsc_data_out_ibuf(12)  (.O (
         image_floue_rsc_data_out_int[12]), .I (image_floue_rsc_data_out[12])) ;
    IBUF \image_floue_rsc_data_out_ibuf(13)  (.O (
         image_floue_rsc_data_out_int[13]), .I (image_floue_rsc_data_out[13])) ;
    IBUF \image_floue_rsc_data_out_ibuf(14)  (.O (
         image_floue_rsc_data_out_int[14]), .I (image_floue_rsc_data_out[14])) ;
    IBUF \image_floue_rsc_data_out_ibuf(15)  (.O (
         image_floue_rsc_data_out_int[15]), .I (image_floue_rsc_data_out[15])) ;
    IBUF \image_floue_rsc_data_out_ibuf(16)  (.O (
         image_floue_rsc_data_out_int[16]), .I (image_floue_rsc_data_out[16])) ;
    IBUF \image_floue_rsc_data_out_ibuf(17)  (.O (
         image_floue_rsc_data_out_int[17]), .I (image_floue_rsc_data_out[17])) ;
    IBUF \image_floue_rsc_data_out_ibuf(18)  (.O (
         image_floue_rsc_data_out_int[18]), .I (image_floue_rsc_data_out[18])) ;
    IBUF \image_floue_rsc_data_out_ibuf(19)  (.O (
         image_floue_rsc_data_out_int[19]), .I (image_floue_rsc_data_out[19])) ;
    IBUF \image_floue_rsc_data_out_ibuf(20)  (.O (
         image_floue_rsc_data_out_int[20]), .I (image_floue_rsc_data_out[20])) ;
    IBUF \image_floue_rsc_data_out_ibuf(21)  (.O (
         image_floue_rsc_data_out_int[21]), .I (image_floue_rsc_data_out[21])) ;
    IBUF \image_floue_rsc_data_out_ibuf(22)  (.O (
         image_floue_rsc_data_out_int[22]), .I (image_floue_rsc_data_out[22])) ;
    IBUF \image_floue_rsc_data_out_ibuf(23)  (.O (
         image_floue_rsc_data_out_int[23]), .I (image_floue_rsc_data_out[23])) ;
    IBUF \image_floue_rsc_data_out_ibuf(24)  (.O (
         image_floue_rsc_data_out_int[24]), .I (image_floue_rsc_data_out[24])) ;
    IBUF \image_floue_rsc_data_out_ibuf(25)  (.O (
         image_floue_rsc_data_out_int[25]), .I (image_floue_rsc_data_out[25])) ;
    IBUF \image_floue_rsc_data_out_ibuf(26)  (.O (
         image_floue_rsc_data_out_int[26]), .I (image_floue_rsc_data_out[26])) ;
    IBUF \image_floue_rsc_data_out_ibuf(27)  (.O (
         image_floue_rsc_data_out_int[27]), .I (image_floue_rsc_data_out[27])) ;
    IBUF \image_floue_rsc_data_out_ibuf(28)  (.O (
         image_floue_rsc_data_out_int[28]), .I (image_floue_rsc_data_out[28])) ;
    IBUF \image_floue_rsc_data_out_ibuf(29)  (.O (
         image_floue_rsc_data_out_int[29]), .I (image_floue_rsc_data_out[29])) ;
    IBUF \image_floue_rsc_data_out_ibuf(30)  (.O (
         image_floue_rsc_data_out_int[30]), .I (image_floue_rsc_data_out[30])) ;
    IBUF \image_floue_rsc_data_out_ibuf(31)  (.O (
         image_floue_rsc_data_out_int[31]), .I (image_floue_rsc_data_out[31])) ;
    IBUF \image_net_rsc_data_out_ibuf(0)  (.O (image_net_rsc_data_out_int[0]), .I (
         image_net_rsc_data_out[0])) ;
    IBUF \image_net_rsc_data_out_ibuf(1)  (.O (image_net_rsc_data_out_int[1]), .I (
         image_net_rsc_data_out[1])) ;
    IBUF \image_net_rsc_data_out_ibuf(2)  (.O (image_net_rsc_data_out_int[2]), .I (
         image_net_rsc_data_out[2])) ;
    IBUF \image_net_rsc_data_out_ibuf(3)  (.O (image_net_rsc_data_out_int[3]), .I (
         image_net_rsc_data_out[3])) ;
    IBUF \image_net_rsc_data_out_ibuf(4)  (.O (image_net_rsc_data_out_int[4]), .I (
         image_net_rsc_data_out[4])) ;
    IBUF \image_net_rsc_data_out_ibuf(5)  (.O (image_net_rsc_data_out_int[5]), .I (
         image_net_rsc_data_out[5])) ;
    IBUF \image_net_rsc_data_out_ibuf(6)  (.O (image_net_rsc_data_out_int[6]), .I (
         image_net_rsc_data_out[6])) ;
    IBUF \image_net_rsc_data_out_ibuf(7)  (.O (image_net_rsc_data_out_int[7]), .I (
         image_net_rsc_data_out[7])) ;
    IBUF \image_net_rsc_data_out_ibuf(8)  (.O (image_net_rsc_data_out_int[8]), .I (
         image_net_rsc_data_out[8])) ;
    IBUF \image_net_rsc_data_out_ibuf(9)  (.O (image_net_rsc_data_out_int[9]), .I (
         image_net_rsc_data_out[9])) ;
    IBUF \image_net_rsc_data_out_ibuf(10)  (.O (image_net_rsc_data_out_int[10])
         , .I (image_net_rsc_data_out[10])) ;
    IBUF \image_net_rsc_data_out_ibuf(11)  (.O (image_net_rsc_data_out_int[11])
         , .I (image_net_rsc_data_out[11])) ;
    IBUF \image_net_rsc_data_out_ibuf(12)  (.O (image_net_rsc_data_out_int[12])
         , .I (image_net_rsc_data_out[12])) ;
    IBUF \image_net_rsc_data_out_ibuf(13)  (.O (image_net_rsc_data_out_int[13])
         , .I (image_net_rsc_data_out[13])) ;
    IBUF \image_net_rsc_data_out_ibuf(14)  (.O (image_net_rsc_data_out_int[14])
         , .I (image_net_rsc_data_out[14])) ;
    IBUF \image_net_rsc_data_out_ibuf(15)  (.O (image_net_rsc_data_out_int[15])
         , .I (image_net_rsc_data_out[15])) ;
    IBUF \image_net_rsc_data_out_ibuf(16)  (.O (image_net_rsc_data_out_int[16])
         , .I (image_net_rsc_data_out[16])) ;
    IBUF \image_net_rsc_data_out_ibuf(17)  (.O (image_net_rsc_data_out_int[17])
         , .I (image_net_rsc_data_out[17])) ;
    IBUF \image_net_rsc_data_out_ibuf(18)  (.O (image_net_rsc_data_out_int[18])
         , .I (image_net_rsc_data_out[18])) ;
    IBUF \image_net_rsc_data_out_ibuf(19)  (.O (image_net_rsc_data_out_int[19])
         , .I (image_net_rsc_data_out[19])) ;
    IBUF \image_net_rsc_data_out_ibuf(20)  (.O (image_net_rsc_data_out_int[20])
         , .I (image_net_rsc_data_out[20])) ;
    IBUF \image_net_rsc_data_out_ibuf(21)  (.O (image_net_rsc_data_out_int[21])
         , .I (image_net_rsc_data_out[21])) ;
    IBUF \image_net_rsc_data_out_ibuf(22)  (.O (image_net_rsc_data_out_int[22])
         , .I (image_net_rsc_data_out[22])) ;
    IBUF \image_net_rsc_data_out_ibuf(23)  (.O (image_net_rsc_data_out_int[23])
         , .I (image_net_rsc_data_out[23])) ;
    IBUF \image_net_rsc_data_out_ibuf(24)  (.O (image_net_rsc_data_out_int[24])
         , .I (image_net_rsc_data_out[24])) ;
    IBUF \image_net_rsc_data_out_ibuf(25)  (.O (image_net_rsc_data_out_int[25])
         , .I (image_net_rsc_data_out[25])) ;
    IBUF \image_net_rsc_data_out_ibuf(26)  (.O (image_net_rsc_data_out_int[26])
         , .I (image_net_rsc_data_out[26])) ;
    IBUF \image_net_rsc_data_out_ibuf(27)  (.O (image_net_rsc_data_out_int[27])
         , .I (image_net_rsc_data_out[27])) ;
    IBUF \image_net_rsc_data_out_ibuf(28)  (.O (image_net_rsc_data_out_int[28])
         , .I (image_net_rsc_data_out[28])) ;
    IBUF \image_net_rsc_data_out_ibuf(29)  (.O (image_net_rsc_data_out_int[29])
         , .I (image_net_rsc_data_out[29])) ;
    IBUF \image_net_rsc_data_out_ibuf(30)  (.O (image_net_rsc_data_out_int[30])
         , .I (image_net_rsc_data_out[30])) ;
    IBUF \image_net_rsc_data_out_ibuf(31)  (.O (image_net_rsc_data_out_int[31])
         , .I (image_net_rsc_data_out[31])) ;
    IBUF rst_ibuf (.O (rst_int), .I (rst)) ;
    INV ix35068z1315 (.O (image_error_rsc_re_1_0), .I (
        \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
    INV ix15434z1315 (.O (depth_rsc_we_1_0), .I (\main_core_inst_fsm_output(10)  
        )) ;
    GND ps_gnd (.G (nx18058z10)) ;
    VCC ps_vcc (.P (nx18058z11)) ;
    main_core_0 main_core_inst (.px1915 (nx60417z1), .px1914 (nx59420z1), .px1913 (
                nx58423z1), .px1912 (nx57426z1), .px1911 (nx56429z1), .px1910 (
                nx55432z1), .px1909 (nx54435z1), .px1908 (nx53438z1), .px1907 (
                nx52441z1), .px1906 (nx51444z1), .px1905 (nx9824z1), .px1904 (
                nx10821z1), .px1903 (nx11818z1), .px1902 (nx12815z1), .px1901 (
                nx13812z1), .px1900 (nx14809z1), .px1899 (nx15806z1), .px1898 (
                nx16803z1), .px1897 (nx17800z1), .px1896 (nx18797z1), .px1895 (
                nx20793z1), .px1894 (nx21790z1), .px1893 (nx22787z1), .px1892 (
                nx23784z1), .px1891 (nx24781z1), .px1890 (nx25778z1), .px1889 (
                nx26775z1), .px1888 (nx27772z1), .px1887 (nx28769z1), .px1886 (
                nx29766z1), .px1885 (nx31762z1), .px1884 (nx32759z1), .px1877 (
                nx51351z1), .px1876 (nx62619z1), .px1875 (nx61622z1), .px1874 (
                nx60625z1), .px1873 (nx59628z1), .px1872 (nx58631z1), .px1871 (
                nx57634z1), .px1870 (nx56637z1), .px1869 (nx55640z1), .px1868 (
                nx54643z1), .px1867 (nx53646z1), .px1866 (nx22882z1), .px1865 (
                nx21885z1), .px1864 (nx20888z1), .px1863 (nx19891z1), .px1862 (
                nx18894z1), .px1861 (nx17897z1), .px1860 (nx16900z1), .px1859 (
                nx19538z1), .px1858 (nx20535z1), .px1857 (nx21532z1), .px1856 (
                nx22529z1), .px1855 (nx23526z1), .px1854 (nx24523z1), .px1853 (
                nx25520z1), .px1852 (nx26517z1), .px1851 (nx27514z1), .px1850 (
                nx28511z1), .px1849 (nx33183z1), .px1848 (nx34180z1), .px1847 (
                nx35177z1), .px1846 (nx36174z1), .px1845 (nx37171z1), .px1844 (
                nx38168z1), .px1843 (nx39165z1), .px1842 (nx40162z1), .px1841 (
                nx41159z1), .px1840 (nx42156z1), .px1839 (nx44152z1), .px1838 (
                nx45149z1), .px1837 (nx46146z1), .px1836 (nx47143z1), .px1835 (
                nx48140z1), .px1834 (nx49137z1), .px1833 (nx50134z1), .px1832 (
                nx51131z1), .px1831 (nx52128z1), .px1830 (nx53125z1), .px1829 (
                nx55121z1), .px1828 (nx56118z1), .px1827 (nx7721z1), .p_nbus_image_error_rsc_data_out_int (
                {image_error_rsc_data_out_int[13],
                image_error_rsc_data_out_int[12],
                image_error_rsc_data_out_int[11],
                image_error_rsc_data_out_int[10],image_error_rsc_data_out_int[9]
                ,image_error_rsc_data_out_int[8],image_error_rsc_data_out_int[7]
                ,image_error_rsc_data_out_int[6],image_error_rsc_data_out_int[5]
                ,image_error_rsc_data_out_int[2],
                image_error_rsc_data_out_int[16],
                image_error_rsc_data_out_int[15],
                image_error_rsc_data_out_int[14],image_error_rsc_data_out_int[4]
                ,image_error_rsc_data_out_int[3],image_error_rsc_data_out_int[1]
                ,image_error_rsc_data_out_int[0],
                image_error_rsc_data_out_int[31],
                image_error_rsc_data_out_int[30],
                image_error_rsc_data_out_int[29],
                image_error_rsc_data_out_int[28],
                image_error_rsc_data_out_int[27],
                image_error_rsc_data_out_int[26],
                image_error_rsc_data_out_int[25],
                image_error_rsc_data_out_int[24],
                image_error_rsc_data_out_int[23],
                image_error_rsc_data_out_int[22],
                image_error_rsc_data_out_int[21],
                image_error_rsc_data_out_int[20],
                image_error_rsc_data_out_int[19],
                image_error_rsc_data_out_int[18],
                image_error_rsc_data_out_int[17]}), .p_nbus_image_net_rsc_data_out_int (
                {image_net_rsc_data_out_int[31],image_net_rsc_data_out_int[30],
                image_net_rsc_data_out_int[29],image_net_rsc_data_out_int[28],
                image_net_rsc_data_out_int[27],image_net_rsc_data_out_int[26],
                image_net_rsc_data_out_int[25],image_net_rsc_data_out_int[24],
                image_net_rsc_data_out_int[23],image_net_rsc_data_out_int[22],
                image_net_rsc_data_out_int[21],image_net_rsc_data_out_int[20],
                image_net_rsc_data_out_int[19],image_net_rsc_data_out_int[18],
                image_net_rsc_data_out_int[17],image_net_rsc_data_out_int[16],
                image_net_rsc_data_out_int[15],image_net_rsc_data_out_int[14],
                image_net_rsc_data_out_int[13],image_net_rsc_data_out_int[12],
                image_net_rsc_data_out_int[11],image_net_rsc_data_out_int[10],
                image_net_rsc_data_out_int[9],image_net_rsc_data_out_int[8],
                image_net_rsc_data_out_int[7],image_net_rsc_data_out_int[6],
                image_net_rsc_data_out_int[5],image_net_rsc_data_out_int[4],
                image_net_rsc_data_out_int[3],image_net_rsc_data_out_int[2],
                image_net_rsc_data_out_int[1],image_net_rsc_data_out_int[0]}), .p_nbus_image_floue_rsc_data_out_int (
                {image_floue_rsc_data_out_int[31],
                image_floue_rsc_data_out_int[30],
                image_floue_rsc_data_out_int[29],
                image_floue_rsc_data_out_int[28],
                image_floue_rsc_data_out_int[27],
                image_floue_rsc_data_out_int[26],
                image_floue_rsc_data_out_int[25],
                image_floue_rsc_data_out_int[24],
                image_floue_rsc_data_out_int[23],
                image_floue_rsc_data_out_int[22],
                image_floue_rsc_data_out_int[21],
                image_floue_rsc_data_out_int[20],
                image_floue_rsc_data_out_int[19],
                image_floue_rsc_data_out_int[18],
                image_floue_rsc_data_out_int[17],
                image_floue_rsc_data_out_int[16],
                image_floue_rsc_data_out_int[15],
                image_floue_rsc_data_out_int[14],
                image_floue_rsc_data_out_int[13],
                image_floue_rsc_data_out_int[12],
                image_floue_rsc_data_out_int[11],
                image_floue_rsc_data_out_int[10],image_floue_rsc_data_out_int[9]
                ,image_floue_rsc_data_out_int[8],image_floue_rsc_data_out_int[7]
                ,image_floue_rsc_data_out_int[6],image_floue_rsc_data_out_int[5]
                ,image_floue_rsc_data_out_int[4],image_floue_rsc_data_out_int[3]
                ,image_floue_rsc_data_out_int[2],image_floue_rsc_data_out_int[1]
                ,image_floue_rsc_data_out_int[0]}), .p_nbus_depth_rsc_addr_1_0 (
                {depth_rsc_addr_1_0[2],depth_rsc_addr_1_0[1],
                depth_rsc_addr_1_0[0]}), .\p_fsm_output(10)   (
                \main_core_inst_fsm_output(10)  ), .p_image_net_rsc_triosy_lz_1_0 (
                image_net_rsc_triosy_lz_1_0), .p_nbus_image_net_rsc_addr_1_0 ({
                image_net_rsc_addr_1_0[0],image_net_rsc_addr_1_0[1],
                image_net_rsc_addr_1_0[2],image_net_rsc_addr_1_0[15],
                image_net_rsc_addr_1_0[14],image_net_rsc_addr_1_0[13],
                image_net_rsc_addr_1_0[12],image_net_rsc_addr_1_0[11],
                image_net_rsc_addr_1_0[10],image_net_rsc_addr_1_0[9],
                image_net_rsc_addr_1_0[8],image_net_rsc_addr_1_0[7],
                image_net_rsc_addr_1_0[6],image_net_rsc_addr_1_0[5],
                image_net_rsc_addr_1_0[4],image_net_rsc_addr_1_0[3]}), .p_rst_int (
                rst_int), .p_clk_int (clk_int), .px1642 (nx18058z1), .px1644 (
                nx18058z2), .px1646 (nx18058z3), .px1648 (nx18058z4), .px1650 (
                nx18058z5), .px1652 (nx18058z6), .px1654 (nx18058z7), .px1656 (
                nx18058z8), .px1658 (nx18058z9), .\p_z_out(8)   (
                \main_core_inst_z_out(8)  ), .\p_z_out(7)   (
                \main_core_inst_z_out(7)  ), .\p_z_out(6)   (
                \main_core_inst_z_out(6)  ), .\p_z_out(5)   (
                \main_core_inst_z_out(5)  ), .\p_z_out(4)   (
                \main_core_inst_z_out(4)  ), .\p_z_out(3)   (
                \main_core_inst_z_out(3)  ), .\p_z_out(2)   (
                \main_core_inst_z_out(2)  ), .\p_z_out(1)   (
                \main_core_inst_z_out(1)  ), .\p_z_out(0)   (
                \main_core_inst_z_out(0)  ), .\p_for_for_mux1h_2_nl(1)   (
                \main_core_inst_for_for_mux1h_2_nl(1)  ), .px1302 (nx18058z10), 
                .px1918 (nx18058z11)) ;
    BUFGP clk_ibuf (.O (clk_int), .I (clk)) ;
    LUT2 ix18058z15973 (.O (nx18058z1), .I0 (\main_core_inst_z_out(8)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15973.INIT = 4'h8;
    LUT2 ix18058z15974 (.O (nx18058z2), .I0 (\main_core_inst_z_out(7)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15974.INIT = 4'h8;
    LUT2 ix18058z15975 (.O (nx18058z3), .I0 (\main_core_inst_z_out(6)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15975.INIT = 4'h8;
    LUT2 ix18058z15976 (.O (nx18058z4), .I0 (\main_core_inst_z_out(5)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15976.INIT = 4'h8;
    LUT2 ix18058z15977 (.O (nx18058z5), .I0 (\main_core_inst_z_out(4)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15977.INIT = 4'h8;
    LUT2 ix18058z15978 (.O (nx18058z6), .I0 (\main_core_inst_z_out(3)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15978.INIT = 4'h8;
    LUT2 ix18058z15979 (.O (nx18058z7), .I0 (\main_core_inst_z_out(2)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15979.INIT = 4'h8;
    LUT2 ix18058z15980 (.O (nx18058z8), .I0 (\main_core_inst_z_out(1)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15980.INIT = 4'h8;
    LUT2 ix18058z15981 (.O (nx18058z9), .I0 (\main_core_inst_z_out(0)  ), .I1 (
         \main_core_inst_for_for_mux1h_2_nl(1)  )) ;
         defparam ix18058z15981.INIT = 4'h8;
endmodule


module main_core_0 ( px1915, px1914, px1913, px1912, px1911, px1910, px1909, 
                     px1908, px1907, px1906, px1905, px1904, px1903, px1902, 
                     px1901, px1900, px1899, px1898, px1897, px1896, px1895, 
                     px1894, px1893, px1892, px1891, px1890, px1889, px1888, 
                     px1887, px1886, px1885, px1884, px1877, px1876, px1875, 
                     px1874, px1873, px1872, px1871, px1870, px1869, px1868, 
                     px1867, px1866, px1865, px1864, px1863, px1862, px1861, 
                     px1860, px1859, px1858, px1857, px1856, px1855, px1854, 
                     px1853, px1852, px1851, px1850, px1849, px1848, px1847, 
                     px1846, px1845, px1844, px1843, px1842, px1841, px1840, 
                     px1839, px1838, px1837, px1836, px1835, px1834, px1833, 
                     px1832, px1831, px1830, px1829, px1828, px1827, 
                     p_nbus_image_error_rsc_data_out_int, 
                     p_nbus_image_net_rsc_data_out_int, 
                     p_nbus_image_floue_rsc_data_out_int, 
                     p_nbus_depth_rsc_addr_1_0, \p_fsm_output(10)  , 
                     p_image_net_rsc_triosy_lz_1_0, 
                     p_nbus_image_net_rsc_addr_1_0, p_rst_int, p_clk_int, px1642, 
                     px1644, px1646, px1648, px1650, px1652, px1654, px1656, 
                     px1658, \p_z_out(8)  , \p_z_out(7)  , \p_z_out(6)  , 
                     \p_z_out(5)  , \p_z_out(4)  , \p_z_out(3)  , \p_z_out(2)  , 
                     \p_z_out(1)  , \p_z_out(0)  , \p_for_for_mux1h_2_nl(1)  , 
                     px1302, px1918 ) ;

    output px1915 ;
    output px1914 ;
    output px1913 ;
    output px1912 ;
    output px1911 ;
    output px1910 ;
    output px1909 ;
    output px1908 ;
    output px1907 ;
    output px1906 ;
    output px1905 ;
    output px1904 ;
    output px1903 ;
    output px1902 ;
    output px1901 ;
    output px1900 ;
    output px1899 ;
    output px1898 ;
    output px1897 ;
    output px1896 ;
    output px1895 ;
    output px1894 ;
    output px1893 ;
    output px1892 ;
    output px1891 ;
    output px1890 ;
    output px1889 ;
    output px1888 ;
    output px1887 ;
    output px1886 ;
    output px1885 ;
    output px1884 ;
    output px1877 ;
    output px1876 ;
    output px1875 ;
    output px1874 ;
    output px1873 ;
    output px1872 ;
    output px1871 ;
    output px1870 ;
    output px1869 ;
    output px1868 ;
    output px1867 ;
    output px1866 ;
    output px1865 ;
    output px1864 ;
    output px1863 ;
    output px1862 ;
    output px1861 ;
    output px1860 ;
    output px1859 ;
    output px1858 ;
    output px1857 ;
    output px1856 ;
    output px1855 ;
    output px1854 ;
    output px1853 ;
    output px1852 ;
    output px1851 ;
    output px1850 ;
    output px1849 ;
    output px1848 ;
    output px1847 ;
    output px1846 ;
    output px1845 ;
    output px1844 ;
    output px1843 ;
    output px1842 ;
    output px1841 ;
    output px1840 ;
    output px1839 ;
    output px1838 ;
    output px1837 ;
    output px1836 ;
    output px1835 ;
    output px1834 ;
    output px1833 ;
    output px1832 ;
    output px1831 ;
    output px1830 ;
    output px1829 ;
    output px1828 ;
    output px1827 ;
    input [31:0]p_nbus_image_error_rsc_data_out_int ;
    input [31:0]p_nbus_image_net_rsc_data_out_int ;
    input [31:0]p_nbus_image_floue_rsc_data_out_int ;
    output [2:0]p_nbus_depth_rsc_addr_1_0 ;
    output \p_fsm_output(10)   ;
    output p_image_net_rsc_triosy_lz_1_0 ;
    output [15:0]p_nbus_image_net_rsc_addr_1_0 ;
    input p_rst_int ;
    input p_clk_int ;
    input px1642 ;
    input px1644 ;
    input px1646 ;
    input px1648 ;
    input px1650 ;
    input px1652 ;
    input px1654 ;
    input px1656 ;
    input px1658 ;
    output \p_z_out(8)   ;
    output \p_z_out(7)   ;
    output \p_z_out(6)   ;
    output \p_z_out(5)   ;
    output \p_z_out(4)   ;
    output \p_z_out(3)   ;
    output \p_z_out(2)   ;
    output \p_z_out(1)   ;
    output \p_z_out(0)   ;
    output \p_for_for_mux1h_2_nl(1)   ;
    input px1302 ;
    input px1918 ;

    wire nx34290z3, nx6053z6, nx6053z5, nx6053z4, nx6053z3, nx6053z2, nx12063z4, 
         nx12062z4, nx12061z4, nx12060z4, nx7975z7, nx7974z3, nx7977z7, 
         nx10394z10, nx10394z12, nx10394z14, nx10394z16, nx10394z18, nx10394z20, 
         nx10394z22, nx10394z24, nx10394z26, nx56495z6, nx11516z5, nx21850z3, 
         nx21850z2, nx23844z3, nx24841z4, nx24841z3, nx24841z2, nx25838z4, 
         nx25838z3, nx25838z2, nx26835z2, nx27832z2, nx4228z2, nx3231z2, 
         nx1235z2, nx238z2, nx64777z2, nx63780z2, nx62783z2, nx61786z2, 
         nx60789z2, nx59792z2, nx58795z2, nx57798z2, nx55802z2, nx54805z2, 
         nx53808z2, nx52811z2, nx51814z2, nx50817z2, nx49820z2, nx48823z2, 
         nx47826z2, nx46829z2, nx5781z2, nx4784z2, nx3787z2, nx2790z2, nx1793z2, 
         nx796z2, nx65335z2, nx64338z2, nx63341z2, nx62344z2, nx7977z4, nx7975z4, 
         nx7976z4, nx56495z5, nx8012z4, nx8012z3, nx8012z2, nx29305z2, nx56495z3, 
         nx64941z2, nx58489z2, nx1399z4, nx64941z3, nx1399z2, nx56495z4, 
         nx21269z2, nx22266z2, nx23263z2, nx21269z3, nx11516z6, nx11516z4, 
         nx23844z2, nx11515z4, nx11515z3, nx11514z4, nx11514z3, nx11510z6, 
         nx11510z5, nx52183z3, nx7973z3, nx7975z6, nx7975z3, nx7976z3, nx7977z3, 
         nx29245z1, nx4943z10, nx28248z1, nx4943z9, nx27251z1, nx4943z8, 
         nx26254z1, nx4943z7, nx25257z1, nx4943z6, nx24260z1, nx4943z5, 
         nx23263z1, nx4943z4, nx22266z1, nx4943z3, nx21269z1, nx4943z2, 
         nx25029z1, nx56642z2, nx24032z1, nx57639z2, nx23035z2, nx11510z4, 
         nx22038z1, nx13034z3, nx21041z1, nx12037z2, nx20044z1, nx11040z2, 
         nx19047z1, nx10043z2, nx18050z1, nx9046z2, nx17053z1, nx23035z1, 
         nx8049z2, nx61480z1, nx60483z1, nx1399z3, nx58489z1, nx64941z4, 
         nx57492z1, nx56495z7, nx56495z2, nx56495z1, nx63944z3, nx65061z2, 
         nx522z2, nx1519z2, nx2516z2, nx3513z2, nx4510z2, nx5507z2, nx6504z2, 
         nx7501z2, nx32296z2, nx29305z1, \fsm_output(1)  , nx31299z1, 
         \main_core_core_fsm_inst_fsm_output(3)  , nx32296z1, \fsm_output(4)  , 
         nx33293z1, \fsm_output(5)  , nx34290z1, \fsm_output(6)  , nx35287z1, 
         \fsm_output(8)  , nx37281z1, \fsm_output(9)  , nx38278z1, 
         \fsm_output(11)  , nx7015z1, \fsm_output(12)  , nx8012z1, nx9009z1, 
         \fsm_output(0)  , nx8049z1;
    wire [5:0]main_core_inst_for_1_for_acc_7_psp_1_sva_1;
    wire nx9046z1, nx10043z1, nx11040z1, nx12037z1, nx13034z2, nx40352z1;
    wire [22:0]main_core_inst_reconstruction_error_for_for_c_sva_31_9_2;
    wire nx41349z1, nx42346z1, nx43343z1, nx44340z2, nx45337z1, nx46334z1, 
         nx47331z1, nx48328z1, nx49325z1, nx55707z1, nx54710z1, nx53713z1, 
         nx52716z1, nx51719z1, nx50722z1, nx49725z1, nx48728z1, nx47731z1, 
         nx46734z1, nx44738z1, nx43741z1, nx42744z1, nx44340z1, nx4577z1;
    wire [31:0]main_core_inst_reconstruction_error_for_l_sva_3;
    wire nx5574z1, nx6571z1, nx7568z1, nx8565z1, nx9562z1, nx10559z1, nx11556z1, 
         nx12553z1, nx13550z1, nx59274z1, nx60271z1, nx61268z1, nx62265z1, 
         nx63262z1, nx64259z1, nx65256z1, nx717z1, nx1714z1, nx2711z1, nx4707z1, 
         nx5704z1, nx6701z1, nx7698z1, nx8695z1, nx9692z1, nx10689z1, nx11686z1, 
         nx12683z1, nx13680z1, nx15676z1, nx16673z2, nx16673z1, 
         \for_1_for_acc_6_psp_1_sva(0)  ;
    wire [4:0]main_core_inst_for_1_for_acc_6_psp_1_sva_1;
    wire nx7974z5, nx7975z8, nx7976z5, nx7977z5, nx13034z1, nx63474z2, nx62477z1, 
         nx59486z1, nx63474z1, \for_1_i_7_0_sva_4(4)  , nx65061z1;
    wire [8:0]main_core_inst_for_for_j_8_0_sva_3;
    wire nx522z1, nx1519z1, nx2516z1, nx3513z1, nx4510z1, nx5507z1, nx6504z1, 
         nx7501z1;
    wire [13:0]main_core_inst_for_for_else_acc_itm_2;
    wire nx6053z1, for_for_if_for_for_if_and_itm_1, nx61860z1;
    wire [31:0]main_core_inst_reconstruction_error_rec_error_sva;
    wire nx60863z1, nx59866z1, nx58869z1, nx57872z1, nx56875z1, nx55878z1, 
         nx54881z1, nx53884z1, nx52887z1, nx52591z1, nx51594z1, nx50597z1, 
         nx49600z1, nx48603z1, nx47606z1, nx46609z1, nx45612z1, nx44615z1, 
         nx43618z1, nx41622z1, nx40625z1, nx39628z1, nx38631z1, nx37634z1, 
         nx36637z1, nx35640z1, nx34643z1, nx33646z1, nx32649z1, nx30653z1, 
         nx29656z1, nx62344z1;
    wire [31:0]main_core_inst_reconstruction_error_rec_error_lpi_6;
    wire nx63341z1, nx64338z1, nx65335z1, nx796z1, nx1793z1, nx2790z1, nx3787z1, 
         nx4784z1, nx5781z1, nx46829z1, nx47826z1, nx48823z1, nx49820z1, 
         nx50817z1, nx51814z1, nx52811z1, nx53808z1, nx54805z1, nx55802z1, 
         nx57798z1, nx58795z1, nx59792z1, nx60789z1, nx61786z1, nx62783z1, 
         nx63780z1, nx64777z1, nx238z1, nx1235z1, nx3231z1, nx4228z1, nx26190z1, 
         exit_reconstruction_error_for_for_sva_1, 
         for_1_for_slc_for_1_for_acc_7_itm_1, nx56642z1;
    wire [8:0]main_core_inst_for_1_for_j_8_0_sva_4;
    wire nx57639z1, nx27832z1, nx26835z1, nx25838z1, nx24841z1, nx23844z1, 
         nx22847z1, nx21850z1, nx5387z1, nx4390z1, nx3393z1, nx2396z1, 
         \for_i_7_0_sva_3(3)  , nx1399z1, \for_i_7_0_sva_3(4)  , nx402z1, 
         \for_i_7_0_sva_3(5)  , nx64941z1, \for_i_7_0_sva_3(6)  , nx63944z2, 
         nx63944z1, \for_i_7_0_sva_3(7)  , nx42790z15, nx42790z14, nx42790z13, 
         nx42790z12, nx42790z11, nx42790z10, nx42790z9, nx42790z8, nx42790z7, 
         nx42790z6, nx42790z5, nx42790z4, nx42790z3, nx42790z2, nx42790z1;
    wire [31:31]main_core_inst_z_out;
    wire \z_out(18)  , \z_out(19)  , \z_out(20)  , \z_out(21)  , \z_out(22)  , 
         \z_out(23)  , \z_out(24)  , \z_out(25)  , \z_out(26)  , \z_out(27)  , 
         \z_out(28)  , \z_out(29)  , \z_out(30)  , \z_out(31)  , nx6176z15, 
         nx6176z14, nx6176z13, nx6176z12, nx6176z11, nx6176z10, nx6176z9, 
         nx6176z8, nx6176z7, nx6176z6, nx6176z5, nx6176z4, nx6176z3, nx6176z2, 
         nx6176z1, nx42790z63, nx42790z62, nx42790z61, nx42790z60, nx42790z59, 
         nx42790z58, nx42790z57, nx42790z56, nx42790z55, nx42790z54, nx42790z53, 
         nx42790z52, nx42790z51, nx42790z50, nx42790z49, nx42790z48, nx42790z47, 
         nx42790z46, nx42790z45, nx42790z44, nx42790z43, nx42790z42, nx42790z41, 
         nx42790z40, nx42790z39, nx42790z38, nx42790z37, nx42790z36, nx42790z35, 
         nx42790z34, nx42790z33, nx42790z32, nx42790z31, nx42790z30, nx42790z29, 
         nx42790z28, nx42790z27, nx42790z26, nx42790z25, nx42790z24, nx42790z23, 
         nx42790z22, nx42790z21, nx42790z20, nx42790z19, nx42790z18, nx42790z17, 
         nx42790z16, nx10394z43, nx10394z42, nx10394z41, nx10394z40, nx10394z39, 
         nx10394z38, nx10394z37, nx10394z36, nx10394z35, nx10394z34, nx10394z33, 
         nx10394z32, nx10394z31, nx10394z30, nx10394z29, nx10394z28, nx10394z27, 
         nx10394z25, nx10394z23, nx10394z21, nx10394z19, nx10394z17, nx10394z15, 
         nx10394z13, nx10394z11, nx10394z9, nx10394z8, nx10394z7, nx10394z6, 
         nx10394z5, nx10394z4, nx10394z3, nx10394z2, nx10394z1, nx6176z81, 
         nx6176z80, nx6176z79, nx6176z78, nx6176z77, nx6176z76, nx6176z75, 
         nx6176z74, nx6176z73, nx6176z72, nx6176z71, nx6176z70, nx6176z69, 
         nx6176z68, nx6176z67, nx6176z66, nx6176z65, nx6176z64, nx6176z63, 
         nx6176z62, nx6176z61, nx6176z60, nx6176z59, nx6176z58, nx6176z57, 
         nx6176z56, nx6176z55, nx6176z54, nx6176z53, nx6176z52, nx6176z51, 
         nx6176z50, nx6176z49, nx6176z48, nx6176z47, nx6176z46, nx6176z45, 
         nx6176z44, nx6176z43, nx6176z42, nx6176z41, nx6176z40, nx6176z39, 
         nx6176z38, nx6176z37, nx6176z36, nx6176z35, nx6176z34, \z_out(14)  , 
         \z_out(15)  , \z_out(16)  , nx6176z33, nx6176z32, nx6176z31, nx6176z30, 
         nx6176z29, nx6176z28, nx6176z27, nx6176z26, nx6176z25, nx6176z24, 
         nx6176z23, nx6176z22, nx6176z21, nx6176z20, nx6176z19, nx6176z18, 
         nx6176z17, nx6176z16;
    wire [12:2]main_core_inst_for_for_else_mul_2_nl;
    wire nx41749z1, nx60377z2, nx60377z1, nx60378z2, nx60378z1, nx60379z2, 
         nx60379z1, nx60380z2, nx60380z1, nx60381z2, nx60381z1, nx60382z2, 
         nx60382z1, nx60383z2, nx60383z1, nx60384z2, nx60384z1, nx60385z2, 
         nx60385z1, nx60386z1, \a(9)  , \a(8)  , nx42839z1, \a(7)  , nx42838z1, 
         nx42837z2, \a(6)  , nx42837z1, nx42836z2, \a(5)  , nx42836z1, nx42835z2, 
         \a(4)  , nx42835z1, nx42834z2, \a(3)  , nx42834z1, nx42833z2, \a(2)  , 
         nx42833z1, nx42832z2, \a(1)  , nx42832z1, nx42831z1, \a(0)  , nx23312z2, 
         image_error_mux1h_nl_0n0s3, nx38388z1, nx23312z1, nx23311z2;
    wire [3:0]main_core_inst_image_error_mux_nl;
    wire nx38387z1, nx23311z1, nx23310z2, nx38386z1, nx23310z1, nx23309z2, 
         nx26274z1, nx23309z1, nx33887z2, nx33887z1, nx33888z2;
    wire [8:0]main_core_inst_image_error_mux1h_2_nl_0n0s3;
    wire nx33888z1, nx33889z2, nx33889z1, nx33890z2, nx33890z1, nx33891z2, 
         nx33891z1, nx33892z2, nx33892z1, nx33893z2, nx33893z1, nx33894z2, 
         nx33894z1, nx33895z2, nx33895z1, nx33896z1, nx52183z2, 
         \reconstruction_error_for_acc_3_nl(8)  , nx7977z6, nx7977z2, nx52183z1, 
         nx7976z6, nx7976z2, nx7977z1, nx7975z5, nx7975z2, nx7976z1, nx7974z4, 
         nx7974z2, nx7975z1, nx7973z4, nx7973z2, nx7974z1, nx7972z3, nx7972z2, 
         nx7973z1, nx7971z1, \reconstruction_error_for_acc_3_nl_0n0s2(0)  , 
         nx7972z1, nx45700z2;
    wire [31:0]main_core_inst_z_out_6;
    wire nx34912z1, nx45700z1, nx45701z2, nx33924z1, nx45701z1, nx46689z2, 
         nx33923z1, nx46689z1, nx46690z2, nx33922z1, nx46690z1, nx46691z2, 
         nx33921z1, nx46691z1, nx46692z2, nx33920z1, nx46692z1, nx46693z2, 
         nx33919z1, nx46693z1, nx46694z2, nx33918z1, nx46694z1, nx46695z2, 
         nx33917z1, nx46695z1, nx46696z2, nx33916z1, nx46696z1, nx46697z2, 
         nx33915z1, nx46697z1, nx46698z2, nx32927z1, nx46698z1, nx47686z2, 
         nx32926z1, nx47686z1, nx47687z2, nx32925z1, nx47687z1, nx47688z2, 
         nx32924z1, nx47688z1, nx47689z2, nx32923z1, nx47689z1, nx47690z2, 
         nx32922z1, nx47690z1, nx47691z2, nx32921z1, nx47691z1, nx47692z2, 
         nx32920z1, nx47692z1, nx47693z2, nx32919z1, nx47693z1, nx47694z2, 
         nx32918z1, nx47694z1, nx47695z2, nx17526z1, nx47695z1, nx42635z2, 
         nx17525z1, nx42635z1, nx42636z2, nx17524z1, nx42636z1, nx42637z2, 
         nx17523z1, nx42637z1, nx42638z2, nx17522z1, nx42638z1, nx42639z2, 
         nx17521z1, nx42639z1, nx42640z2, nx17520z1, nx42640z1, nx42641z2, 
         nx17519z1, nx42641z1, nx42642z2, nx17518z1, nx42642z1, nx42643z2, 
         nx17517z1, nx42643z1, nx42644z1, not_fsm_output_8, nx50036z2, 
         \main_core_core_fsm_inst_reconstruction_error_for_C_0_tr0_0n0s3(7)  , 
         nx39524z3, nx39524z2, nx50036z1, nx39523z3, nx39523z2, nx39524z1, 
         nx39522z3, nx39522z2, nx39523z1, nx39521z3, nx39521z2, nx39522z1, 
         nx39520z3, nx39520z2, nx39521z1, nx39519z2, nx39520z1, nx39519z3, 
         nx39519z1, nx34672z3, nx34672z2, nx34290z2, nx35660z3, nx35660z2, 
         nx34672z1, nx35661z3, nx35661z2, nx35660z1, nx35662z3, nx35662z2, 
         nx35661z1, nx35663z3, nx35663z2, nx35662z1, nx35664z3, nx35664z2, 
         nx35663z1, nx35665z3, nx35665z2, nx35664z1, nx35666z3, nx35666z2, 
         nx35665z1, nx35667z3, nx35667z2, nx35666z1, nx35668z3, nx35668z2, 
         nx35667z1, nx35669z3, nx35669z2, nx35668z1, nx36657z3, nx36657z2, 
         nx35669z1, nx36658z3, nx36658z2, nx36657z1, nx36659z3, nx36659z2, 
         nx36658z1, nx36660z3, nx36660z2, nx36659z1, nx36661z3, nx36661z2, 
         nx36660z1, nx36662z3, nx36662z2, nx36661z1, nx36663z3, nx36663z2, 
         nx36662z1, nx36664z3, nx36664z2, nx36663z1, nx36665z3, nx36665z2, 
         nx36664z1, nx36666z3, nx36666z2, nx36665z1, nx12058z3, nx12058z2, 
         nx36666z1, nx12059z3, nx12059z2, nx12058z1, nx12060z3, nx12060z2, 
         nx12059z1, nx12061z3, nx12061z2, nx12060z1, nx12062z3, nx12062z2, 
         nx12061z1, nx12063z3, nx12063z2, nx12062z1, nx12064z3, nx12064z2, 
         nx12063z1, nx12065z3, nx12065z2, nx12064z1, nx12066z3, nx12066z2, 
         nx12065z1, nx12067z2, nx12067z1, nx12066z1;
    wire \z_out(13)  ;
    wire \for_for_else_acc_itm_2_14n1s1(13)  , nx18473z1;
    wire \z_out(12)  ;
    wire \for_for_else_acc_itm_2_14n1s1(12)  , nx18474z1;
    wire \z_out(11)  ;
    wire \for_for_else_acc_itm_2_14n1s1(11)  , nx18475z1;
    wire \z_out(10)  ;
    wire \for_for_else_acc_itm_2_14n1s1(10)  , nx18476z1;
    wire \z_out(9)  ;
    wire \for_for_else_acc_itm_2_14n1s1(9)  , nx42716z1;
    wire [8:0]main_core_inst_for_for_if_acc_nl;
    wire nx42715z1, nx42714z1, nx42713z1, nx42712z1, nx42711z2, nx42711z1, 
         nx42710z2, nx42710z1, nx42709z2, nx42709z1, nx42708z2, nx42708z1, 
         nx42707z1, nx11516z3;
    wire [7:0]main_core_inst_z_out_2;
    wire nx48644z1, nx11516z2, nx11516z1, nx11515z2, nx11515z1, nx11514z2, 
         nx11514z1, nx11513z2, nx11512z2, nx11513z1, nx11512z3, nx11512z1, 
         nx11511z2, nx11510z2, nx11511z1, nx11510z3, nx40591z2, nx40591z1, 
         nx55667z2, nx55667z1, nx55666z2, nx55666z1, nx25634z2, nx25634z1, 
         nx25633z2, nx25633z1, nx25632z2, nx25632z1, nx25631z2, nx25631z1, 
         nx25630z2, nx25629z2, nx25630z1, nx25629z3, nx25628z2, nx25629z1, 
         nx25628z3, nx25627z2, nx25628z1, nx25627z3, nx25626z2, nx25627z1, 
         nx25626z3, nx25625z1, nx25626z1, nx25625z2;
    wire [8:0]main_core_inst_z_out_8;
    wire [22:0]main_core_inst_reconstruction_error_for_for_c_mux_nl;
    wire nx4943z1;
    wire [540:0] \$dummy ;




    inc_32_0 reconstruction_error_for_for_c_mux_nl_inc32_10 (.a ({nx4943z1,
             \$dummy [0],\$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],
             \$dummy [5],\$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],
             \$dummy [10],\$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
             \$dummy [15],\$dummy [16],\$dummy [17],\$dummy [18],\$dummy [19],
             \$dummy [20],\$dummy [21],\$dummy [22],\$dummy [23],\$dummy [24],
             \$dummy [25],\$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29],
             \$dummy [30]}), .d ({
             main_core_inst_reconstruction_error_for_for_c_mux_nl[0],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[1],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[2],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[3],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[4],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[5],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[6],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[7],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[8],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[9],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[10],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[11],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[12],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[13],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[14],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[15],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[16],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[17],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[18],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[19],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[20],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[21],
             main_core_inst_reconstruction_error_for_for_c_mux_nl[22],
             main_core_inst_z_out_8[0],main_core_inst_z_out_8[1],
             main_core_inst_z_out_8[2],main_core_inst_z_out_8[3],
             main_core_inst_z_out_8[4],main_core_inst_z_out_8[5],
             main_core_inst_z_out_8[6],main_core_inst_z_out_8[7],
             main_core_inst_z_out_8[8]}), .\p_reconstruction_error_for_for_c_sva_31_9_2(21)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[1]), .\p_for_for_mux1h_2_nl(1)   (
             \p_for_for_mux1h_2_nl(1)  ), .\p_reconstruction_error_for_l_sva_3(30)   (
             main_core_inst_reconstruction_error_for_l_sva_3[1]), .\p_reconstruction_error_for_for_c_sva_31_9_2(20)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[2]), .\p_reconstruction_error_for_l_sva_3(29)   (
             main_core_inst_reconstruction_error_for_l_sva_3[2]), .\p_reconstruction_error_for_for_c_sva_31_9_2(19)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[3]), .\p_reconstruction_error_for_l_sva_3(28)   (
             main_core_inst_reconstruction_error_for_l_sva_3[3]), .\p_reconstruction_error_for_for_c_sva_31_9_2(18)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[4]), .\p_reconstruction_error_for_l_sva_3(27)   (
             main_core_inst_reconstruction_error_for_l_sva_3[4]), .\p_reconstruction_error_for_for_c_sva_31_9_2(17)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[5]), .\p_reconstruction_error_for_l_sva_3(26)   (
             main_core_inst_reconstruction_error_for_l_sva_3[5]), .\p_reconstruction_error_for_for_c_sva_31_9_2(16)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[6]), .\p_reconstruction_error_for_l_sva_3(25)   (
             main_core_inst_reconstruction_error_for_l_sva_3[6]), .\p_reconstruction_error_for_for_c_sva_31_9_2(15)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[7]), .\p_reconstruction_error_for_l_sva_3(24)   (
             main_core_inst_reconstruction_error_for_l_sva_3[7]), .\p_reconstruction_error_for_for_c_sva_31_9_2(14)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[8]), .\p_reconstruction_error_for_l_sva_3(23)   (
             main_core_inst_reconstruction_error_for_l_sva_3[8]), .\p_reconstruction_error_for_for_c_sva_31_9_2(13)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[9]), .\p_reconstruction_error_for_l_sva_3(22)   (
             main_core_inst_reconstruction_error_for_l_sva_3[9]), .\p_reconstruction_error_for_for_c_sva_31_9_2(12)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[10]), .\p_reconstruction_error_for_l_sva_3(21)   (
             main_core_inst_reconstruction_error_for_l_sva_3[10]), .\p_reconstruction_error_for_for_c_sva_31_9_2(11)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[11]), .\p_reconstruction_error_for_l_sva_3(20)   (
             main_core_inst_reconstruction_error_for_l_sva_3[11]), .\p_reconstruction_error_for_for_c_sva_31_9_2(10)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[12]), .\p_reconstruction_error_for_l_sva_3(19)   (
             main_core_inst_reconstruction_error_for_l_sva_3[12]), .\p_reconstruction_error_for_for_c_sva_31_9_2(9)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[13]), .\p_reconstruction_error_for_l_sva_3(18)   (
             main_core_inst_reconstruction_error_for_l_sva_3[13]), .\p_reconstruction_error_for_for_c_sva_31_9_2(8)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[14]), .\p_reconstruction_error_for_l_sva_3(17)   (
             main_core_inst_reconstruction_error_for_l_sva_3[14]), .\p_reconstruction_error_for_for_c_sva_31_9_2(7)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[15]), .\p_reconstruction_error_for_l_sva_3(16)   (
             main_core_inst_reconstruction_error_for_l_sva_3[15]), .\p_reconstruction_error_for_for_c_sva_31_9_2(6)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[16]), .\p_reconstruction_error_for_l_sva_3(15)   (
             main_core_inst_reconstruction_error_for_l_sva_3[16]), .\p_reconstruction_error_for_for_c_sva_31_9_2(5)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[17]), .\p_reconstruction_error_for_l_sva_3(14)   (
             main_core_inst_reconstruction_error_for_l_sva_3[17]), .\p_reconstruction_error_for_for_c_sva_31_9_2(4)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[18]), .\p_reconstruction_error_for_l_sva_3(13)   (
             main_core_inst_reconstruction_error_for_l_sva_3[18]), .\p_reconstruction_error_for_for_c_sva_31_9_2(3)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[19]), .\p_reconstruction_error_for_l_sva_3(12)   (
             main_core_inst_reconstruction_error_for_l_sva_3[19]), .\p_reconstruction_error_for_for_c_sva_31_9_2(2)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[20]), .\p_reconstruction_error_for_l_sva_3(11)   (
             main_core_inst_reconstruction_error_for_l_sva_3[20]), .\p_reconstruction_error_for_for_c_sva_31_9_2(1)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[21]), .\p_reconstruction_error_for_l_sva_3(10)   (
             main_core_inst_reconstruction_error_for_l_sva_3[21]), .\p_reconstruction_error_for_for_c_sva_31_9_2(0)   (
             main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[22]), .\p_reconstruction_error_for_l_sva_3(9)   (
             main_core_inst_reconstruction_error_for_l_sva_3[22]), .\p_reconstruction_error_for_l_sva_3(8)   (
             main_core_inst_reconstruction_error_for_l_sva_3[23]), .px2488 (
             nx4943z2), .\p_reconstruction_error_for_l_sva_3(7)   (
             main_core_inst_reconstruction_error_for_l_sva_3[24]), .px2489 (
             nx4943z3), .\p_reconstruction_error_for_l_sva_3(6)   (
             main_core_inst_reconstruction_error_for_l_sva_3[25]), .px2490 (
             nx4943z4), .\p_reconstruction_error_for_l_sva_3(5)   (
             main_core_inst_reconstruction_error_for_l_sva_3[26]), .px2491 (
             nx4943z5), .\p_reconstruction_error_for_l_sva_3(4)   (
             main_core_inst_reconstruction_error_for_l_sva_3[27]), .px2492 (
             nx4943z6), .\p_reconstruction_error_for_l_sva_3(3)   (
             main_core_inst_reconstruction_error_for_l_sva_3[28]), .px2493 (
             nx4943z7), .\p_reconstruction_error_for_l_sva_3(2)   (
             main_core_inst_reconstruction_error_for_l_sva_3[29]), .px2494 (
             nx4943z8), .\p_reconstruction_error_for_l_sva_3(1)   (
             main_core_inst_reconstruction_error_for_l_sva_3[30]), .px2495 (
             nx4943z9), .\p_reconstruction_error_for_l_sva_3(0)   (
             main_core_inst_reconstruction_error_for_l_sva_3[31]), .px2496 (
             nx4943z10)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_0 (.O (
          p_nbus_image_net_rsc_addr_1_0[0]), .CI (px1302), .LI (nx25625z2)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_1 (.O (
          p_nbus_image_net_rsc_addr_1_0[1]), .CI (nx25626z1), .LI (nx25626z3)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_2 (.O (
          p_nbus_image_net_rsc_addr_1_0[2]), .CI (nx25627z1), .LI (nx25627z3)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_3 (.O (
          p_nbus_image_net_rsc_addr_1_0[3]), .CI (nx25628z1), .LI (nx25628z3)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_4 (.O (
          p_nbus_image_net_rsc_addr_1_0[4]), .CI (nx25629z1), .LI (nx25629z3)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_5 (.O (
          p_nbus_image_net_rsc_addr_1_0[5]), .CI (nx25630z1), .LI (nx25630z2)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_6 (.O (
          p_nbus_image_net_rsc_addr_1_0[6]), .CI (nx25631z1), .LI (nx25631z2)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_7 (.O (
          p_nbus_image_net_rsc_addr_1_0[7]), .CI (nx25632z1), .LI (nx25632z2)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_8 (.O (
          p_nbus_image_net_rsc_addr_1_0[8]), .CI (nx25633z1), .LI (nx25633z2)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_9 (.O (
          p_nbus_image_net_rsc_addr_1_0[9]), .CI (nx25634z1), .LI (nx25634z2)) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_10 (.O (
          p_nbus_image_net_rsc_addr_1_0[10]), .CI (nx55666z1), .LI (nx55666z2)
          ) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_11 (.O (
          p_nbus_image_net_rsc_addr_1_0[11]), .CI (nx55667z1), .LI (nx55667z2)
          ) ;
    XORCY image_net_rsci_addr_d_add13_4_xorcy_12 (.O (
          p_nbus_image_net_rsc_addr_1_0[12]), .CI (nx40591z1), .LI (nx40591z2)
          ) ;
    XORCY z_out_2_add8_5_xorcy_0 (.O (main_core_inst_z_out_2[0]), .CI (px1302), 
          .LI (nx11510z3)) ;
    XORCY z_out_2_add8_5_xorcy_1 (.O (main_core_inst_z_out_2[1]), .CI (nx11511z1
          ), .LI (nx11511z2)) ;
    XORCY z_out_2_add8_5_xorcy_2 (.O (main_core_inst_z_out_2[2]), .CI (nx11512z1
          ), .LI (nx11512z3)) ;
    XORCY z_out_2_add8_5_xorcy_3 (.O (main_core_inst_z_out_2[3]), .CI (nx11513z1
          ), .LI (nx11513z2)) ;
    XORCY z_out_2_add8_5_xorcy_4 (.O (main_core_inst_z_out_2[4]), .CI (nx11514z1
          ), .LI (nx11514z2)) ;
    XORCY z_out_2_add8_5_xorcy_5 (.O (main_core_inst_z_out_2[5]), .CI (nx11515z1
          ), .LI (nx11515z2)) ;
    XORCY z_out_2_add8_5_xorcy_6 (.O (main_core_inst_z_out_2[6]), .CI (nx11516z1
          ), .LI (nx11516z2)) ;
    XORCY z_out_2_add8_5_xorcy_7 (.O (main_core_inst_z_out_2[7]), .CI (nx48644z1
          ), .LI (nx11516z3)) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_0 (.O (
          main_core_inst_for_for_if_acc_nl[0]), .CI (px1302), .LI (nx42707z1)) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_1 (.O (
          main_core_inst_for_for_if_acc_nl[1]), .CI (nx42708z1), .LI (nx42708z2)
          ) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_2 (.O (
          main_core_inst_for_for_if_acc_nl[2]), .CI (nx42709z1), .LI (nx42709z2)
          ) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_3 (.O (
          main_core_inst_for_for_if_acc_nl[3]), .CI (nx42710z1), .LI (nx42710z2)
          ) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_4 (.O (
          main_core_inst_for_for_if_acc_nl[4]), .CI (nx42711z1), .LI (nx42711z2)
          ) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_5 (.O (
          main_core_inst_for_for_if_acc_nl[5]), .CI (nx42712z1), .LI (
          \p_z_out(5)  )) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_6 (.O (
          main_core_inst_for_for_if_acc_nl[6]), .CI (nx42713z1), .LI (
          \p_z_out(6)  )) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_7 (.O (
          main_core_inst_for_for_if_acc_nl[7]), .CI (nx42714z1), .LI (
          \p_z_out(7)  )) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_8 (.O (
          main_core_inst_for_for_if_acc_nl[8]), .CI (nx42715z1), .LI (
          \p_z_out(8)  )) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_9 (.O (
          \for_for_else_acc_itm_2_14n1s1(9)  ), .CI (nx42716z1), .LI (\z_out(9)  
          )) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_10 (.O (
          \for_for_else_acc_itm_2_14n1s1(10)  ), .CI (nx18476z1), .LI (
          \z_out(10)  )) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_11 (.O (
          \for_for_else_acc_itm_2_14n1s1(11)  ), .CI (nx18475z1), .LI (
          \z_out(11)  )) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_12 (.O (
          \for_for_else_acc_itm_2_14n1s1(12)  ), .CI (nx18474z1), .LI (
          \z_out(12)  )) ;
    XORCY for_for_else_acc_itm_2_add14_14i1_xorcy_13 (.O (
          \for_for_else_acc_itm_2_14n1s1(13)  ), .CI (nx18473z1), .LI (
          \z_out(13)  )) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_30 (.O (nx34290z2), .CI (
          nx34672z1), .DI (nx34672z2), .S (nx34672z3)) ;
    GND ps_gnd (.G (nx39519z1)) ;
    VCC ps_vcc (.P (nx39519z3)) ;
    XORCY xorcy_0_9 (.O (
          \main_core_core_fsm_inst_reconstruction_error_for_C_0_tr0_0n0s3(7)  )
          , .CI (nx50036z1), .LI (nx50036z2)) ;
    XORCY z_out_6_add33_6_xorcy_0 (.O (main_core_inst_z_out_6[0]), .CI (
          not_fsm_output_8), .LI (nx42644z1)) ;
    XORCY z_out_6_add33_6_xorcy_1 (.O (main_core_inst_z_out_6[1]), .CI (
          nx42643z1), .LI (nx42643z2)) ;
    XORCY z_out_6_add33_6_xorcy_2 (.O (main_core_inst_z_out_6[2]), .CI (
          nx42642z1), .LI (nx42642z2)) ;
    XORCY z_out_6_add33_6_xorcy_3 (.O (main_core_inst_z_out_6[3]), .CI (
          nx42641z1), .LI (nx42641z2)) ;
    XORCY z_out_6_add33_6_xorcy_4 (.O (main_core_inst_z_out_6[4]), .CI (
          nx42640z1), .LI (nx42640z2)) ;
    XORCY z_out_6_add33_6_xorcy_5 (.O (main_core_inst_z_out_6[5]), .CI (
          nx42639z1), .LI (nx42639z2)) ;
    XORCY z_out_6_add33_6_xorcy_6 (.O (main_core_inst_z_out_6[6]), .CI (
          nx42638z1), .LI (nx42638z2)) ;
    XORCY z_out_6_add33_6_xorcy_7 (.O (main_core_inst_z_out_6[7]), .CI (
          nx42637z1), .LI (nx42637z2)) ;
    XORCY z_out_6_add33_6_xorcy_8 (.O (main_core_inst_z_out_6[8]), .CI (
          nx42636z1), .LI (nx42636z2)) ;
    XORCY z_out_6_add33_6_xorcy_9 (.O (main_core_inst_z_out_6[9]), .CI (
          nx42635z1), .LI (nx42635z2)) ;
    XORCY z_out_6_add33_6_xorcy_10 (.O (main_core_inst_z_out_6[10]), .CI (
          nx47695z1), .LI (nx47695z2)) ;
    XORCY z_out_6_add33_6_xorcy_11 (.O (main_core_inst_z_out_6[11]), .CI (
          nx47694z1), .LI (nx47694z2)) ;
    XORCY z_out_6_add33_6_xorcy_12 (.O (main_core_inst_z_out_6[12]), .CI (
          nx47693z1), .LI (nx47693z2)) ;
    XORCY z_out_6_add33_6_xorcy_13 (.O (main_core_inst_z_out_6[13]), .CI (
          nx47692z1), .LI (nx47692z2)) ;
    XORCY z_out_6_add33_6_xorcy_14 (.O (main_core_inst_z_out_6[14]), .CI (
          nx47691z1), .LI (nx47691z2)) ;
    XORCY z_out_6_add33_6_xorcy_15 (.O (main_core_inst_z_out_6[15]), .CI (
          nx47690z1), .LI (nx47690z2)) ;
    XORCY z_out_6_add33_6_xorcy_16 (.O (main_core_inst_z_out_6[16]), .CI (
          nx47689z1), .LI (nx47689z2)) ;
    XORCY z_out_6_add33_6_xorcy_17 (.O (main_core_inst_z_out_6[17]), .CI (
          nx47688z1), .LI (nx47688z2)) ;
    XORCY z_out_6_add33_6_xorcy_18 (.O (main_core_inst_z_out_6[18]), .CI (
          nx47687z1), .LI (nx47687z2)) ;
    XORCY z_out_6_add33_6_xorcy_19 (.O (main_core_inst_z_out_6[19]), .CI (
          nx47686z1), .LI (nx47686z2)) ;
    XORCY z_out_6_add33_6_xorcy_20 (.O (main_core_inst_z_out_6[20]), .CI (
          nx46698z1), .LI (nx46698z2)) ;
    XORCY z_out_6_add33_6_xorcy_21 (.O (main_core_inst_z_out_6[21]), .CI (
          nx46697z1), .LI (nx46697z2)) ;
    XORCY z_out_6_add33_6_xorcy_22 (.O (main_core_inst_z_out_6[22]), .CI (
          nx46696z1), .LI (nx46696z2)) ;
    XORCY z_out_6_add33_6_xorcy_23 (.O (main_core_inst_z_out_6[23]), .CI (
          nx46695z1), .LI (nx46695z2)) ;
    XORCY z_out_6_add33_6_xorcy_24 (.O (main_core_inst_z_out_6[24]), .CI (
          nx46694z1), .LI (nx46694z2)) ;
    XORCY z_out_6_add33_6_xorcy_25 (.O (main_core_inst_z_out_6[25]), .CI (
          nx46693z1), .LI (nx46693z2)) ;
    XORCY z_out_6_add33_6_xorcy_26 (.O (main_core_inst_z_out_6[26]), .CI (
          nx46692z1), .LI (nx46692z2)) ;
    XORCY z_out_6_add33_6_xorcy_27 (.O (main_core_inst_z_out_6[27]), .CI (
          nx46691z1), .LI (nx46691z2)) ;
    XORCY z_out_6_add33_6_xorcy_28 (.O (main_core_inst_z_out_6[28]), .CI (
          nx46690z1), .LI (nx46690z2)) ;
    XORCY z_out_6_add33_6_xorcy_29 (.O (main_core_inst_z_out_6[29]), .CI (
          nx46689z1), .LI (nx46689z2)) ;
    XORCY z_out_6_add33_6_xorcy_30 (.O (main_core_inst_z_out_6[30]), .CI (
          nx45701z1), .LI (nx45701z2)) ;
    XORCY z_out_6_add33_6_xorcy_31 (.O (main_core_inst_z_out_6[31]), .CI (
          nx45700z1), .LI (nx45700z2)) ;
    XORCY reconstruction_error_for_acc_3_nl_add9_1_xorcy_7 (.O (
          \reconstruction_error_for_acc_3_nl(8)  ), .CI (nx52183z1), .LI (
          nx52183z2)) ;
    XORCY modgen_add_4_xorcy_0 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[0]), .CI (px1302), .LI (
          nx33896z1)) ;
    XORCY modgen_add_4_xorcy_1 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[1]), .CI (nx33895z1), .LI (
          nx33895z2)) ;
    XORCY modgen_add_4_xorcy_2 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[2]), .CI (nx33894z1), .LI (
          nx33894z2)) ;
    XORCY modgen_add_4_xorcy_3 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[3]), .CI (nx33893z1), .LI (
          nx33893z2)) ;
    XORCY modgen_add_4_xorcy_4 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[4]), .CI (nx33892z1), .LI (
          nx33892z2)) ;
    XORCY modgen_add_4_xorcy_5 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[5]), .CI (nx33891z1), .LI (
          nx33891z2)) ;
    XORCY modgen_add_4_xorcy_6 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[6]), .CI (nx33890z1), .LI (
          nx33890z2)) ;
    XORCY modgen_add_4_xorcy_7 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[7]), .CI (nx33889z1), .LI (
          nx33889z2)) ;
    XORCY modgen_add_4_xorcy_8 (.O (
          main_core_inst_image_error_mux1h_2_nl_0n0s3[8]), .CI (nx33888z1), .LI (
          nx33888z2)) ;
    XORCY modgen_add_4_xorcy_9 (.O (main_core_inst_image_error_mux_nl[0]), .CI (
          nx33887z1), .LI (nx33887z2)) ;
    XORCY modgen_add_4_xorcy_10 (.O (main_core_inst_image_error_mux_nl[1]), .CI (
          nx23309z1), .LI (nx23309z2)) ;
    XORCY modgen_add_4_xorcy_11 (.O (main_core_inst_image_error_mux_nl[2]), .CI (
          nx23310z1), .LI (nx23310z2)) ;
    XORCY modgen_add_4_xorcy_12 (.O (main_core_inst_image_error_mux_nl[3]), .CI (
          nx23311z1), .LI (nx23311z2)) ;
    XORCY modgen_add_4_xorcy_13 (.O (image_error_mux1h_nl_0n0s3), .CI (nx23312z1
          ), .LI (nx23312z2)) ;
    XORCY ix456_xorcy_0 (.O (\a(0)  ), .CI (px1302), .LI (nx42831z1)) ;
    XORCY ix456_xorcy_1 (.O (\a(1)  ), .CI (nx42832z1), .LI (nx42832z2)) ;
    XORCY ix456_xorcy_2 (.O (\a(2)  ), .CI (nx42833z1), .LI (nx42833z2)) ;
    XORCY ix456_xorcy_3 (.O (\a(3)  ), .CI (nx42834z1), .LI (nx42834z2)) ;
    XORCY ix456_xorcy_4 (.O (\a(4)  ), .CI (nx42835z1), .LI (nx42835z2)) ;
    XORCY ix456_xorcy_5 (.O (\a(5)  ), .CI (nx42836z1), .LI (nx42836z2)) ;
    XORCY ix456_xorcy_6 (.O (\a(6)  ), .CI (nx42837z1), .LI (nx42837z2)) ;
    XORCY ix456_xorcy_7 (.O (\a(7)  ), .CI (nx42838z1), .LI (
          main_core_inst_for_for_j_8_0_sva_3[5])) ;
    XORCY ix456_xorcy_8 (.O (\a(8)  ), .CI (nx42839z1), .LI (
          main_core_inst_for_for_j_8_0_sva_3[6])) ;
    MUXCY ix456_muxcy_8 (.O (\a(9)  ), .CI (nx42839z1), .DI (px1302), .S (
          main_core_inst_for_for_j_8_0_sva_3[6])) ;
    XORCY ix486_xorcy_0 (.O (main_core_inst_for_for_else_mul_2_nl[2]), .CI (
          px1302), .LI (nx60386z1)) ;
    XORCY ix486_xorcy_1 (.O (main_core_inst_for_for_else_mul_2_nl[3]), .CI (
          nx60385z1), .LI (nx60385z2)) ;
    XORCY ix486_xorcy_2 (.O (main_core_inst_for_for_else_mul_2_nl[4]), .CI (
          nx60384z1), .LI (nx60384z2)) ;
    XORCY ix486_xorcy_3 (.O (main_core_inst_for_for_else_mul_2_nl[5]), .CI (
          nx60383z1), .LI (nx60383z2)) ;
    XORCY ix486_xorcy_4 (.O (main_core_inst_for_for_else_mul_2_nl[6]), .CI (
          nx60382z1), .LI (nx60382z2)) ;
    XORCY ix486_xorcy_5 (.O (main_core_inst_for_for_else_mul_2_nl[7]), .CI (
          nx60381z1), .LI (nx60381z2)) ;
    XORCY ix486_xorcy_6 (.O (main_core_inst_for_for_else_mul_2_nl[8]), .CI (
          nx60380z1), .LI (nx60380z2)) ;
    XORCY ix486_xorcy_7 (.O (main_core_inst_for_for_else_mul_2_nl[9]), .CI (
          nx60379z1), .LI (nx60379z2)) ;
    XORCY ix486_xorcy_8 (.O (main_core_inst_for_for_else_mul_2_nl[10]), .CI (
          nx60378z1), .LI (nx60378z2)) ;
    XORCY ix486_xorcy_9 (.O (main_core_inst_for_for_else_mul_2_nl[11]), .CI (
          nx60377z1), .LI (nx60377z2)) ;
    XORCY ix486_xorcy_10 (.O (main_core_inst_for_for_else_mul_2_nl[12]), .CI (
          nx41749z1), .LI (\a(8)  )) ;
    FDRE \reg_for_i_7_0_sva_3(7)  (.Q (\for_i_7_0_sva_3(7)  ), .C (p_clk_int), .CE (
         nx63944z1), .D (nx63944z2), .R (p_rst_int)) ;
    FDRE \reg_for_i_7_0_sva_3(6)  (.Q (\for_i_7_0_sva_3(6)  ), .C (p_clk_int), .CE (
         nx63944z1), .D (nx64941z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_7_0_sva_3(5)  (.Q (\for_i_7_0_sva_3(5)  ), .C (p_clk_int), .CE (
         nx63944z1), .D (nx402z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_7_0_sva_3(4)  (.Q (\for_i_7_0_sva_3(4)  ), .C (p_clk_int), .CE (
         nx63944z1), .D (nx1399z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_7_0_sva_3(3)  (.Q (\for_i_7_0_sva_3(3)  ), .C (p_clk_int), .CE (
         nx63944z1), .D (nx2396z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_7_0_sva_3(2)  (.Q (p_nbus_image_net_rsc_addr_1_0[13]), .C (
         p_clk_int), .CE (nx63944z1), .D (nx3393z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_7_0_sva_3(1)  (.Q (p_nbus_image_net_rsc_addr_1_0[14]), .C (
         p_clk_int), .CE (nx63944z1), .D (nx4390z1), .R (p_rst_int)) ;
    FDRE \reg_for_i_7_0_sva_3(0)  (.Q (p_nbus_image_net_rsc_addr_1_0[15]), .C (
         p_clk_int), .CE (nx63944z1), .D (nx5387z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_i_7_0_sva_4(4)  (.Q (\for_1_i_7_0_sva_4(4)  ), .C (p_clk_int
         ), .CE (nx63474z1), .D (nx59486z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_i_7_0_sva_4(1)  (.Q (p_nbus_depth_rsc_addr_1_0[1]), .C (
         p_clk_int), .CE (nx63474z1), .D (nx62477z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_i_7_0_sva_4(0)  (.Q (p_nbus_depth_rsc_addr_1_0[0]), .C (
         p_clk_int), .CE (nx63474z1), .D (nx63474z2), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_6_psp_1_sva_1(4)  (.Q (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[0]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx7977z5), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_6_psp_1_sva_1(3)  (.Q (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[1]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx7976z5), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_6_psp_1_sva_1(2)  (.Q (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[2]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx7975z8), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_6_psp_1_sva_1(1)  (.Q (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[3]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx7974z5), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_6_psp_1_sva_1(0)  (.Q (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[4]), .C (p_clk_int), .CE (
         nx13034z1), .D (\for_1_for_acc_6_psp_1_sva(0)  ), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(31)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[0]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx16673z2), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(30)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[1]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx15676z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(29)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[2]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx13680z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(28)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[3]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx12683z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(27)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[4]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx11686z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(26)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[5]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx10689z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(25)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[6]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx9692z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(24)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[7]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx8695z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(23)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[8]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx7698z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(22)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[9]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx6701z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(21)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[10]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx5704z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(20)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[11]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx4707z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(19)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[12]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx2711z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(18)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[13]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx1714z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(17)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[14]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx717z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(16)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[15]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx65256z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(15)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[16]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx64259z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(14)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[17]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx63262z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(13)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[18]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx62265z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(12)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[19]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx61268z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(11)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[20]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx60271z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(10)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[21]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx59274z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(9)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[22]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx13550z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(8)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[23]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx12553z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(7)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[24]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx11556z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(6)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[25]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx10559z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(5)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[26]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx9562z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(4)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[27]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx8565z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(3)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[28]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx7568z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(2)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[29]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx6571z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(1)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[30]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx5574z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_l_sva_3(0)  (.Q (
         main_core_inst_reconstruction_error_for_l_sva_3[31]), .C (p_clk_int), .CE (
         nx16673z1), .D (nx4577z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(22)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[0]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx42744z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(21)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[1]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx43741z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(20)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[2]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx44738z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(19)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[3]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx46734z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(18)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[4]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx47731z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(17)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[5]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx48728z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(16)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[6]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx49725z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(15)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[7]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx50722z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(14)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[8]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx51719z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(13)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[9]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx52716z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(12)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[10]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx53713z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(11)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[11]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx54710z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(10)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[12]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx55707z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(9)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[13]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx49325z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(8)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[14]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx48328z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(7)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[15]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx47331z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(6)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[16]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx46334z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(5)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[17]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx45337z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(4)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[18]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx44340z2), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(3)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[19]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx43343z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(2)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[20]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx42346z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(1)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[21]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx41349z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_31_9_2(0)  (.Q (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[22]), .C (
         p_clk_int), .CE (nx44340z1), .D (nx40352z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_7_psp_1_sva_1(0)  (.Q (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx13034z2), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_7_psp_1_sva_1(1)  (.Q (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx12037z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_7_psp_1_sva_1(2)  (.Q (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx11040z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_7_psp_1_sva_1(3)  (.Q (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[3]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx10043z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_7_psp_1_sva_1(4)  (.Q (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[4]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx9046z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_acc_7_psp_1_sva_1(5)  (.Q (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[5]), .C (p_clk_int), .CE (
         nx13034z1), .D (nx8049z1), .R (p_rst_int)) ;
    FDRE reg_for_for_slc_for_for_acc_7_itm (.Q (nx32296z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (main_core_inst_z_out_2[7]), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(8)  (.Q (nx7501z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx21850z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(7)  (.Q (nx6504z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx22847z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(6)  (.Q (nx5507z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx23844z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(5)  (.Q (nx4510z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx24841z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(4)  (.Q (nx3513z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx25838z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(3)  (.Q (nx2516z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx26835z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(2)  (.Q (nx1519z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx27832z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(1)  (.Q (nx522z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx57639z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_4(0)  (.Q (nx65061z2), .C (p_clk_int), .CE (
         \fsm_output(1)  ), .D (nx56642z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(8)  (.Q (nx8049z2), .C (p_clk_int), .CE (
         nx23035z1), .D (nx17053z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(7)  (.Q (nx9046z2), .C (p_clk_int), .CE (
         nx23035z1), .D (nx18050z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(6)  (.Q (nx10043z2), .C (p_clk_int), .CE (
         nx23035z1), .D (nx19047z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(5)  (.Q (nx11040z2), .C (p_clk_int), .CE (
         nx23035z1), .D (nx20044z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(4)  (.Q (nx12037z2), .C (p_clk_int), .CE (
         nx23035z1), .D (nx21041z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(3)  (.Q (nx13034z3), .C (p_clk_int), .CE (
         nx23035z1), .D (nx22038z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(2)  (.Q (nx11510z4), .C (p_clk_int), .CE (
         nx23035z1), .D (nx23035z2), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(1)  (.Q (nx57639z2), .C (p_clk_int), .CE (
         nx23035z1), .D (nx24032z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva(0)  (.Q (nx56642z2), .C (p_clk_int), .CE (
         nx23035z1), .D (nx25029z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(8)  (.Q (nx4943z2), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx21269z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(7)  (.Q (nx4943z3), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx22266z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(6)  (.Q (nx4943z4), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx23263z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(5)  (.Q (nx4943z5), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx24260z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(4)  (.Q (nx4943z6), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx25257z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(3)  (.Q (nx4943z7), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx26254z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(2)  (.Q (nx4943z8), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx27251z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(1)  (.Q (nx4943z9), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx28248z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_for_for_c_sva_8_0_2(0)  (.Q (nx4943z10), .C (
         p_clk_int), .CE (not_fsm_output_8), .D (nx29245z1), .R (p_rst_int)) ;
    LUT6 ix52183z1312 (.O (nx52183z2), .I0 (nx7977z3), .I1 (nx7976z3), .I2 (
         nx7975z3), .I3 (nx7975z6), .I4 (nx7973z3), .I5 (nx52183z3)) ;
         defparam ix52183z1312.INIT = 64'hFFFFFFFFFFFFFFFE;
    LUT5 ix25625z49975 (.O (nx25625z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \for_i_7_0_sva_3(3)  ), .I2 (main_core_inst_for_for_j_8_0_sva_3[8]), .I3 (
         \p_z_out(0)  ), .I4 (nx1399z3)) ;
         defparam ix25625z49975.INIT = 32'h14BEBE14;
    LUT5 ix25626z49975 (.O (nx25626z3), .I0 (\p_fsm_output(10)  ), .I1 (
         \for_i_7_0_sva_3(4)  ), .I2 (main_core_inst_for_for_j_8_0_sva_3[7]), .I3 (
         \for_1_i_7_0_sva_4(4)  ), .I4 (\p_z_out(1)  )) ;
         defparam ix25626z49975.INIT = 32'h14BEBE14;
    LUT5 ix25627z46855 (.O (nx25627z3), .I0 (\p_fsm_output(10)  ), .I1 (
         \for_i_7_0_sva_3(5)  ), .I2 (\p_z_out(2)  ), .I3 (
         main_core_inst_for_for_else_mul_2_nl[2]), .I4 (nx64941z4)) ;
         defparam ix25627z46855.INIT = 32'h1B4EB1E4;
    LUT5 ix25628z46855 (.O (nx25628z3), .I0 (\p_fsm_output(10)  ), .I1 (
         \for_i_7_0_sva_3(6)  ), .I2 (\p_z_out(3)  ), .I3 (
         main_core_inst_for_for_else_mul_2_nl[3]), .I4 (nx56495z7)) ;
         defparam ix25628z46855.INIT = 32'h1B4EB1E4;
    LUT5 ix25629z46855 (.O (nx25629z3), .I0 (\p_fsm_output(10)  ), .I1 (
         \for_i_7_0_sva_3(7)  ), .I2 (\p_z_out(4)  ), .I3 (
         main_core_inst_for_for_else_mul_2_nl[4]), .I4 (nx63944z3)) ;
         defparam ix25629z46855.INIT = 32'h1B4EB1E4;
    LUT6 ix11510z23058 (.O (nx11510z3), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (\p_for_for_mux1h_2_nl(1)  ), .I3 (nx11510z4), .I4 (
         nx11510z5), .I5 (nx11510z6)) ;
         defparam ix11510z23058.INIT = 64'h1001FE45100154EF;
    LUT5 ix11511z803 (.O (nx11511z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (main_core_inst_for_1_for_acc_7_psp_1_sva_1[0])
         , .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (nx26835z1)) ;
         defparam ix11511z803.INIT = 32'h10EFFE01;
    LUT5 ix11512z974 (.O (nx11512z3), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (main_core_inst_for_1_for_acc_7_psp_1_sva_1[1])
         , .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (nx25838z1)) ;
         defparam ix11512z974.INIT = 32'h1045FEAB;
    LUT5 ix11513z803 (.O (nx11513z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (main_core_inst_for_1_for_acc_7_psp_1_sva_1[2])
         , .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (nx24841z1)) ;
         defparam ix11513z803.INIT = 32'h10EFFE01;
    LUT6 ix11514z49101 (.O (nx11514z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (main_core_inst_for_1_for_acc_7_psp_1_sva_1[3])
         , .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (nx11514z3), .I5 (nx11514z4)) ;
         defparam ix11514z49101.INIT = 64'h1001FEEF1001BAAB;
    LUT6 ix11515z5411 (.O (nx11515z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (main_core_inst_for_1_for_acc_7_psp_1_sva_1[4])
         , .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (nx11515z3), .I5 (nx11515z4)) ;
         defparam ix11515z5411.INIT = 64'hFEEFBAAB54451001;
    LUT6 ix11516z52971 (.O (nx11516z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[5]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (nx11516z3), .I3 (nx23844z2), .I4 (
         nx11516z4), .I5 (nx11516z6)) ;
         defparam ix11516z52971.INIT = 64'h393939C93939C9C9;
    LUT2 ix42707z1320 (.O (nx42707z1), .I0 (\p_z_out(0)  ), .I1 (
         \for_i_7_0_sva_3(3)  )) ;
         defparam ix42707z1320.INIT = 4'h6;
    LUT2 ix42708z1320 (.O (nx42708z2), .I0 (\p_z_out(1)  ), .I1 (
         \for_i_7_0_sva_3(4)  )) ;
         defparam ix42708z1320.INIT = 4'h6;
    LUT2 ix42709z1320 (.O (nx42709z2), .I0 (\p_z_out(2)  ), .I1 (
         \for_i_7_0_sva_3(5)  )) ;
         defparam ix42709z1320.INIT = 4'h6;
    LUT2 ix42710z1320 (.O (nx42710z2), .I0 (\p_z_out(3)  ), .I1 (
         \for_i_7_0_sva_3(6)  )) ;
         defparam ix42710z1320.INIT = 4'h6;
    LUT2 ix42711z1320 (.O (nx42711z2), .I0 (\p_z_out(4)  ), .I1 (
         \for_i_7_0_sva_3(7)  )) ;
         defparam ix42711z1320.INIT = 4'h6;
    LUT6 ix12067z1279 (.O (nx12067z2), .I0 (p_nbus_depth_rsc_addr_1_0[0]), .I1 (
         \p_fsm_output(10)  ), .I2 (\fsm_output(9)  ), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx56642z2), .I5 (nx12067z1)) ;
         defparam ix12067z1279.INIT = 64'h23230023DCDCFFDC;
    LUT5 ix12066z18967 (.O (nx12066z3), .I0 (p_nbus_depth_rsc_addr_1_0[1]), .I1 (
         \fsm_output(9)  ), .I2 (\p_for_for_mux1h_2_nl(1)  ), .I3 (nx57639z2), .I4 (
         nx12066z2)) ;
         defparam ix12066z18967.INIT = 32'hBB0B44F4;
    LUT5 ix12059z25713 (.O (nx12059z3), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(9)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[23]), .I3 (
         main_core_inst_z_out_2[6]), .I4 (main_core_inst_z_out_8[0])) ;
         defparam ix12059z25713.INIT = 32'h0A1B5F4E;
    LUT3 ix12058z1354 (.O (nx12058z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[22]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[22])) ;
         defparam ix12058z1354.INIT = 8'h27;
    LUT3 ix36666z1354 (.O (nx36666z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[21]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[21])) ;
         defparam ix36666z1354.INIT = 8'h27;
    LUT3 ix36665z1354 (.O (nx36665z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[20]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[20])) ;
         defparam ix36665z1354.INIT = 8'h27;
    LUT3 ix36664z1354 (.O (nx36664z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[19]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[19])) ;
         defparam ix36664z1354.INIT = 8'h27;
    LUT3 ix36663z1354 (.O (nx36663z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[18]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[18])) ;
         defparam ix36663z1354.INIT = 8'h27;
    LUT3 ix36662z1354 (.O (nx36662z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[17]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[17])) ;
         defparam ix36662z1354.INIT = 8'h27;
    LUT3 ix36661z1354 (.O (nx36661z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[16]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[16])) ;
         defparam ix36661z1354.INIT = 8'h27;
    LUT3 ix36660z1354 (.O (nx36660z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[15]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[15])) ;
         defparam ix36660z1354.INIT = 8'h27;
    LUT3 ix36659z1354 (.O (nx36659z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[14]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[14])) ;
         defparam ix36659z1354.INIT = 8'h27;
    LUT3 ix36658z1354 (.O (nx36658z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[13]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[13])) ;
         defparam ix36658z1354.INIT = 8'h27;
    LUT3 ix36657z1354 (.O (nx36657z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[12]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[12])) ;
         defparam ix36657z1354.INIT = 8'h27;
    LUT3 ix35669z1354 (.O (nx35669z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[11]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[11])) ;
         defparam ix35669z1354.INIT = 8'h27;
    LUT3 ix35668z1354 (.O (nx35668z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[10]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[10])) ;
         defparam ix35668z1354.INIT = 8'h27;
    LUT3 ix35667z1354 (.O (nx35667z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[9]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[9])) ;
         defparam ix35667z1354.INIT = 8'h27;
    LUT3 ix35666z1354 (.O (nx35666z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[8]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[8])) ;
         defparam ix35666z1354.INIT = 8'h27;
    LUT3 ix35665z1354 (.O (nx35665z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[7]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[7])) ;
         defparam ix35665z1354.INIT = 8'h27;
    LUT3 ix35664z1354 (.O (nx35664z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[6]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[6])) ;
         defparam ix35664z1354.INIT = 8'h27;
    LUT3 ix35663z1354 (.O (nx35663z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[5]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[5])) ;
         defparam ix35663z1354.INIT = 8'h27;
    LUT3 ix35662z1354 (.O (nx35662z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[4]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[4])) ;
         defparam ix35662z1354.INIT = 8'h27;
    LUT3 ix35661z1354 (.O (nx35661z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[3]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[3])) ;
         defparam ix35661z1354.INIT = 8'h27;
    LUT3 ix35660z1354 (.O (nx35660z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[2]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[2])) ;
         defparam ix35660z1354.INIT = 8'h27;
    LUT3 ix34672z1354 (.O (nx34672z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[1]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[1])) ;
         defparam ix34672z1354.INIT = 8'h27;
    LUT5 ix42644z59217 (.O (nx42644z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[31]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[0]), .I3 (
         p_nbus_image_net_rsc_data_out_int[0]), .I4 (\p_z_out(0)  )) ;
         defparam ix42644z59217.INIT = 32'hD11DE22E;
    LUT5 ix42643z59216 (.O (nx42643z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[30]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[1]), .I3 (
         p_nbus_image_net_rsc_data_out_int[1]), .I4 (\p_z_out(1)  )) ;
         defparam ix42643z59216.INIT = 32'hD11DE22E;
    LUT5 ix42642z59216 (.O (nx42642z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[29]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[2]), .I3 (
         p_nbus_image_net_rsc_data_out_int[2]), .I4 (\p_z_out(2)  )) ;
         defparam ix42642z59216.INIT = 32'hD11DE22E;
    LUT5 ix42641z59216 (.O (nx42641z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[28]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[3]), .I3 (
         p_nbus_image_net_rsc_data_out_int[3]), .I4 (\p_z_out(3)  )) ;
         defparam ix42641z59216.INIT = 32'hD11DE22E;
    LUT5 ix42640z59216 (.O (nx42640z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[27]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[4]), .I3 (
         p_nbus_image_net_rsc_data_out_int[4]), .I4 (\p_z_out(4)  )) ;
         defparam ix42640z59216.INIT = 32'hD11DE22E;
    LUT5 ix42639z59216 (.O (nx42639z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[26]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[5]), .I3 (
         p_nbus_image_net_rsc_data_out_int[5]), .I4 (\p_z_out(5)  )) ;
         defparam ix42639z59216.INIT = 32'hD11DE22E;
    LUT5 ix42638z59216 (.O (nx42638z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[25]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[6]), .I3 (
         p_nbus_image_net_rsc_data_out_int[6]), .I4 (\p_z_out(6)  )) ;
         defparam ix42638z59216.INIT = 32'hD11DE22E;
    LUT5 ix42637z59216 (.O (nx42637z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[24]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[7]), .I3 (
         p_nbus_image_net_rsc_data_out_int[7]), .I4 (\p_z_out(7)  )) ;
         defparam ix42637z59216.INIT = 32'hD11DE22E;
    LUT5 ix42636z59216 (.O (nx42636z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[23]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[8]), .I3 (
         p_nbus_image_net_rsc_data_out_int[8]), .I4 (\p_z_out(8)  )) ;
         defparam ix42636z59216.INIT = 32'hD11DE22E;
    LUT5 ix42635z59216 (.O (nx42635z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[22]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[9]), .I3 (
         p_nbus_image_net_rsc_data_out_int[9]), .I4 (\z_out(9)  )) ;
         defparam ix42635z59216.INIT = 32'hD11DE22E;
    LUT5 ix47695z59216 (.O (nx47695z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[21]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[10]), .I3 (
         p_nbus_image_net_rsc_data_out_int[10]), .I4 (\z_out(10)  )) ;
         defparam ix47695z59216.INIT = 32'hD11DE22E;
    LUT5 ix47694z59216 (.O (nx47694z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[20]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[11]), .I3 (
         p_nbus_image_net_rsc_data_out_int[11]), .I4 (\z_out(11)  )) ;
         defparam ix47694z59216.INIT = 32'hD11DE22E;
    LUT5 ix47693z59216 (.O (nx47693z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[19]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[12]), .I3 (
         p_nbus_image_net_rsc_data_out_int[12]), .I4 (\z_out(12)  )) ;
         defparam ix47693z59216.INIT = 32'hD11DE22E;
    LUT5 ix47692z59216 (.O (nx47692z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[18]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[13]), .I3 (
         p_nbus_image_net_rsc_data_out_int[13]), .I4 (\z_out(13)  )) ;
         defparam ix47692z59216.INIT = 32'hD11DE22E;
    LUT5 ix47691z59216 (.O (nx47691z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[17]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[14]), .I3 (
         p_nbus_image_net_rsc_data_out_int[14]), .I4 (\z_out(14)  )) ;
         defparam ix47691z59216.INIT = 32'hD11DE22E;
    LUT5 ix47690z59216 (.O (nx47690z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[16]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[15]), .I3 (
         p_nbus_image_net_rsc_data_out_int[15]), .I4 (\z_out(15)  )) ;
         defparam ix47690z59216.INIT = 32'hD11DE22E;
    LUT5 ix47689z59216 (.O (nx47689z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[15]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[16]), .I3 (
         p_nbus_image_net_rsc_data_out_int[16]), .I4 (\z_out(16)  )) ;
         defparam ix47689z59216.INIT = 32'hD11DE22E;
    LUT5 ix47688z59216 (.O (nx47688z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[14]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[17]), .I3 (
         p_nbus_image_net_rsc_data_out_int[17]), .I4 (main_core_inst_z_out[31])
         ) ;
         defparam ix47688z59216.INIT = 32'hD11DE22E;
    LUT5 ix47687z59216 (.O (nx47687z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[13]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[18]), .I3 (
         p_nbus_image_net_rsc_data_out_int[18]), .I4 (\z_out(18)  )) ;
         defparam ix47687z59216.INIT = 32'hD11DE22E;
    LUT5 ix47686z59216 (.O (nx47686z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[12]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[19]), .I3 (
         p_nbus_image_net_rsc_data_out_int[19]), .I4 (\z_out(19)  )) ;
         defparam ix47686z59216.INIT = 32'hD11DE22E;
    LUT5 ix46698z59216 (.O (nx46698z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[11]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[20]), .I3 (
         p_nbus_image_net_rsc_data_out_int[20]), .I4 (\z_out(20)  )) ;
         defparam ix46698z59216.INIT = 32'hD11DE22E;
    LUT5 ix46697z59216 (.O (nx46697z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[10]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[21]), .I3 (
         p_nbus_image_net_rsc_data_out_int[21]), .I4 (\z_out(21)  )) ;
         defparam ix46697z59216.INIT = 32'hD11DE22E;
    LUT5 ix46696z59216 (.O (nx46696z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[9]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[22]), .I3 (
         p_nbus_image_net_rsc_data_out_int[22]), .I4 (\z_out(22)  )) ;
         defparam ix46696z59216.INIT = 32'hD11DE22E;
    LUT5 ix46695z59216 (.O (nx46695z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[8]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[23]), .I3 (
         p_nbus_image_net_rsc_data_out_int[23]), .I4 (\z_out(23)  )) ;
         defparam ix46695z59216.INIT = 32'hD11DE22E;
    LUT5 ix46694z59216 (.O (nx46694z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[7]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[24]), .I3 (
         p_nbus_image_net_rsc_data_out_int[24]), .I4 (\z_out(24)  )) ;
         defparam ix46694z59216.INIT = 32'hD11DE22E;
    LUT5 ix46693z59216 (.O (nx46693z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[6]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[25]), .I3 (
         p_nbus_image_net_rsc_data_out_int[25]), .I4 (\z_out(25)  )) ;
         defparam ix46693z59216.INIT = 32'hD11DE22E;
    LUT5 ix46692z59216 (.O (nx46692z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[5]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[26]), .I3 (
         p_nbus_image_net_rsc_data_out_int[26]), .I4 (\z_out(26)  )) ;
         defparam ix46692z59216.INIT = 32'hD11DE22E;
    LUT5 ix46691z59216 (.O (nx46691z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[4]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[27]), .I3 (
         p_nbus_image_net_rsc_data_out_int[27]), .I4 (\z_out(27)  )) ;
         defparam ix46691z59216.INIT = 32'hD11DE22E;
    LUT5 ix46690z59216 (.O (nx46690z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[3]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[28]), .I3 (
         p_nbus_image_net_rsc_data_out_int[28]), .I4 (\z_out(28)  )) ;
         defparam ix46690z59216.INIT = 32'hD11DE22E;
    LUT5 ix46689z59216 (.O (nx46689z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[2]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[29]), .I3 (
         p_nbus_image_net_rsc_data_out_int[29]), .I4 (\z_out(29)  )) ;
         defparam ix46689z59216.INIT = 32'hD11DE22E;
    LUT5 ix45701z59216 (.O (nx45701z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[1]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[30]), .I3 (
         p_nbus_image_net_rsc_data_out_int[30]), .I4 (\z_out(30)  )) ;
         defparam ix45701z59216.INIT = 32'hD11DE22E;
    LUT5 ix45700z59216 (.O (nx45700z2), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[0]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[31]), .I3 (
         p_nbus_image_net_rsc_data_out_int[31]), .I4 (\z_out(31)  )) ;
         defparam ix45700z59216.INIT = 32'hD11DE22E;
    LUT3 ix7973z1466 (.O (nx7973z4), .I0 (nx1399z3), .I1 (nx7972z2), .I2 (
         nx7973z3)) ;
         defparam ix7973z1466.INIT = 8'h96;
    LUT2 ix42831z1320 (.O (nx42831z1), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[0]), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[8])) ;
         defparam ix42831z1320.INIT = 4'h6;
    LUT2 ix42832z1320 (.O (nx42832z2), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[1]), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[7])) ;
         defparam ix42832z1320.INIT = 4'h6;
    LUT2 ix42833z1320 (.O (nx42833z2), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[2]), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[0])) ;
         defparam ix42833z1320.INIT = 4'h6;
    LUT2 ix42834z1320 (.O (nx42834z2), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[1])) ;
         defparam ix42834z1320.INIT = 4'h6;
    LUT2 ix42835z1320 (.O (nx42835z2), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[2])) ;
         defparam ix42835z1320.INIT = 4'h6;
    LUT2 ix42836z1320 (.O (nx42836z2), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3])) ;
         defparam ix42836z1320.INIT = 4'h6;
    LUT2 ix42837z1320 (.O (nx42837z2), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[6]), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[4])) ;
         defparam ix42837z1320.INIT = 4'h6;
    LUT2 ix60386z1320 (.O (nx60386z1), .I0 (\a(0)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[8])) ;
         defparam ix60386z1320.INIT = 4'h6;
    LUT2 ix60385z1320 (.O (nx60385z2), .I0 (\a(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[7])) ;
         defparam ix60385z1320.INIT = 4'h6;
    LUT2 ix60384z1320 (.O (nx60384z2), .I0 (\a(2)  ), .I1 (\a(0)  )) ;
         defparam ix60384z1320.INIT = 4'h6;
    LUT2 ix60383z1320 (.O (nx60383z2), .I0 (\a(3)  ), .I1 (\a(1)  )) ;
         defparam ix60383z1320.INIT = 4'h6;
    LUT2 ix60382z1320 (.O (nx60382z2), .I0 (\a(4)  ), .I1 (\a(2)  )) ;
         defparam ix60382z1320.INIT = 4'h6;
    LUT2 ix60381z1320 (.O (nx60381z2), .I0 (\a(5)  ), .I1 (\a(3)  )) ;
         defparam ix60381z1320.INIT = 4'h6;
    LUT2 ix60380z1320 (.O (nx60380z2), .I0 (\a(6)  ), .I1 (\a(4)  )) ;
         defparam ix60380z1320.INIT = 4'h6;
    LUT2 ix60379z1320 (.O (nx60379z2), .I0 (\a(7)  ), .I1 (\a(5)  )) ;
         defparam ix60379z1320.INIT = 4'h6;
    LUT2 ix60378z1320 (.O (nx60378z2), .I0 (\a(8)  ), .I1 (\a(6)  )) ;
         defparam ix60378z1320.INIT = 4'h6;
    LUT2 ix60377z1320 (.O (nx60377z2), .I0 (\a(9)  ), .I1 (\a(7)  )) ;
         defparam ix60377z1320.INIT = 4'h6;
    INV ix30615z1315 (.O (\for_1_for_acc_6_psp_1_sva(0)  ), .I (nx1399z3)) ;
    INV ix7971z1315 (.O (\reconstruction_error_for_acc_3_nl_0n0s2(0)  ), .I (
        p_nbus_depth_rsc_addr_1_0[0])) ;
    INV ix42644z1315 (.O (not_fsm_output_8), .I (\fsm_output(8)  )) ;
    INV ix13034z1316 (.O (nx13034z2), .I (nx13034z3)) ;
    (* HLUTNM = "LUT62_1_41" *)
    LUT5 ix52183z23331 (.O (nx52183z3), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \fsm_output(5)  ), .I4 (main_core_inst_for_for_j_8_0_sva_3[1])) ;
         defparam ix52183z23331.INIT = 32'h56FF5600;
    (* HLUTNM = "LUT62_1_48" *)
    LUT3 ix29245z1491 (.O (nx29245z1), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         nx56642z2), .I2 (main_core_inst_z_out_8[8])) ;
         defparam ix29245z1491.INIT = 8'hB1;
    (* HLUTNM = "LUT62_1_48" *)
    LUT4 ix28248z48557 (.O (nx28248z1), .I0 (main_core_inst_z_out_8[7]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (nx57639z2), .I3 (nx56642z2)) ;
         defparam ix28248z48557.INIT = 16'hB88B;
    (* HLUTNM = "LUT62_1_38" *)
    LUT5 ix27251z37082 (.O (nx27251z1), .I0 (main_core_inst_z_out_8[6]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (nx11510z4), .I3 (nx57639z2), .I4 (
         nx56642z2)) ;
         defparam ix27251z37082.INIT = 32'h8B8B8BB8;
    LUT6 ix26254z51943 (.O (nx26254z1), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I1 (
         main_core_inst_z_out_8[5]), .I2 (\p_for_for_mux1h_2_nl(1)  ), .I3 (
         nx11510z4), .I4 (nx57639z2), .I5 (nx56642z2)) ;
         defparam ix26254z51943.INIT = 64'hCAC5CAC5CAC5C5C5;
    LUT5 ix25257z62907 (.O (nx25257z1), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I2 (
         main_core_inst_z_out_8[4]), .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (
         nx21269z3)) ;
         defparam ix25257z62907.INIT = 32'hF0AAF099;
    LUT6 ix24260z44747 (.O (nx24260z1), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I3 (
         main_core_inst_z_out_8[3]), .I4 (\p_for_for_mux1h_2_nl(1)  ), .I5 (
         nx21269z3)) ;
         defparam ix24260z44747.INIT = 64'hFF00AAAAFF00A9A9;
    LUT6 ix23263z45004 (.O (nx23263z1), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[3]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2]), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I3 (
         main_core_inst_z_out_8[2]), .I4 (\p_for_for_mux1h_2_nl(1)  ), .I5 (
         nx23263z2)) ;
         defparam ix23263z45004.INIT = 64'hFF00A9A9FF00AAAA;
    LUT4 ix22266z37082 (.O (nx22266z1), .I0 (main_core_inst_z_out_8[1]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[4]), .I3 (nx22266z2)) ;
         defparam ix22266z37082.INIT = 16'h8BB8;
    LUT4 ix21269z37082 (.O (nx21269z1), .I0 (main_core_inst_z_out_8[0]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[5]), .I3 (nx21269z2)) ;
         defparam ix21269z37082.INIT = 16'h8BB8;
    (* HLUTNM = "LUT62_1_90" *)
    LUT2 ix25029z1322 (.O (nx25029z1), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[8])) ;
         defparam ix25029z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_99" *)
    LUT2 ix24032z1322 (.O (nx24032z1), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[7])) ;
         defparam ix24032z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_88" *)
    LUT2 ix23035z1323 (.O (nx23035z2), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[6])) ;
         defparam ix23035z1323.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_98" *)
    LUT2 ix22038z1322 (.O (nx22038z1), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[5])) ;
         defparam ix22038z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_87" *)
    LUT2 ix21041z1322 (.O (nx21041z1), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[4])) ;
         defparam ix21041z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_87" *)
    LUT2 ix20044z1322 (.O (nx20044z1), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[3])) ;
         defparam ix20044z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_88" *)
    LUT2 ix19047z1322 (.O (nx19047z1), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[2])) ;
         defparam ix19047z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_90" *)
    LUT2 ix18050z1322 (.O (nx18050z1), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[1])) ;
         defparam ix18050z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_89" *)
    LUT2 ix17053z1322 (.O (nx17053z1), .I0 (\fsm_output(11)  ), .I1 (
         main_core_inst_for_1_for_j_8_0_sva_4[0])) ;
         defparam ix17053z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_34" *)
    LUT3 ix23035z1568 (.O (nx23035z1), .I0 (\fsm_output(12)  ), .I1 (
         \fsm_output(11)  ), .I2 (\fsm_output(4)  )) ;
         defparam ix23035z1568.INIT = 8'hFE;
    (* HLUTNM = "LUT62_1_24" *)
    LUT4 ix61480z9522 (.O (nx61480z1), .I0 (nx56495z4), .I1 (p_rst_int), .I2 (
         \fsm_output(12)  ), .I3 (p_nbus_depth_rsc_addr_1_0[2])) ;
         defparam ix61480z9522.INIT = 16'h2010;
    LUT6 ix58489z2342 (.O (nx58489z1), .I0 (p_rst_int), .I1 (\fsm_output(12)  )
         , .I2 (nx64941z3), .I3 (nx1399z4), .I4 (nx56495z4), .I5 (nx58489z2)) ;
         defparam ix58489z2342.INIT = 64'h0404044004040404;
    (* HLUTNM = "LUT62_1_49" *)
    LUT3 ix57492z1330 (.O (nx57492z1), .I0 (nx64941z2), .I1 (p_rst_int), .I2 (
         \fsm_output(12)  )) ;
         defparam ix57492z1330.INIT = 8'h10;
    (* HLUTNM = "LUT62_1_49" *)
    LUT4 ix56495z5443 (.O (nx56495z2), .I0 (nx56495z3), .I1 (p_rst_int), .I2 (
         \fsm_output(12)  ), .I3 (nx63944z3)) ;
         defparam ix56495z5443.INIT = 16'h1020;
    (* HLUTNM = "LUT62_1_45" *)
    LUT3 ix56495z1568 (.O (nx56495z1), .I0 (p_rst_int), .I1 (\fsm_output(12)  )
         , .I2 (\fsm_output(4)  )) ;
         defparam ix56495z1568.INIT = 8'hFE;
    (* HLUTNM = "LUT62_1_42" *)
    LUT5 ix29305z494 (.O (nx29305z1), .I0 (\fsm_output(4)  ), .I1 (
         \fsm_output(0)  ), .I2 (\main_core_core_fsm_inst_fsm_output(3)  ), .I3 (
         nx32296z2), .I4 (nx29305z2)) ;
         defparam ix29305z494.INIT = 32'hFEEEFCCC;
    (* HLUTNM = "LUT62_1_102" *)
    LUT2 ix32296z1316 (.O (nx32296z1), .I0 (
         \main_core_core_fsm_inst_fsm_output(3)  ), .I1 (nx32296z2)) ;
         defparam ix32296z1316.INIT = 4'h2;
    (* HLUTNM = "LUT62_1_34" *)
    LUT5 ix33293z530 (.O (nx33293z1), .I0 (\fsm_output(12)  ), .I1 (
         \fsm_output(11)  ), .I2 (\fsm_output(4)  ), .I3 (
         for_1_for_slc_for_1_for_acc_7_itm_1), .I4 (nx29305z2)) ;
         defparam ix33293z530.INIT = 32'hEEAAFCF0;
    (* HLUTNM = "LUT62_1_29" *)
    LUT4 ix35287z54060 (.O (nx35287z1), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(6)  ), .I2 (exit_reconstruction_error_for_for_sva_1), .I3 (
         \main_core_core_fsm_inst_reconstruction_error_for_C_0_tr0_0n0s3(7)  )
         ) ;
         defparam ix35287z54060.INIT = 16'hCE0A;
    (* HLUTNM = "LUT62_1_29" *)
    LUT4 ix37281z42510 (.O (nx37281z1), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(6)  ), .I2 (exit_reconstruction_error_for_for_sva_1), .I3 (
         \main_core_core_fsm_inst_reconstruction_error_for_C_0_tr0_0n0s3(7)  )
         ) ;
         defparam ix37281z42510.INIT = 16'hA0EC;
    (* HLUTNM = "LUT62_1_89" *)
    LUT2 ix7015z1316 (.O (nx7015z1), .I0 (\fsm_output(11)  ), .I1 (
         for_1_for_slc_for_1_for_acc_7_itm_1)) ;
         defparam ix7015z1316.INIT = 4'h2;
    LUT6 ix8012z1444 (.O (nx8012z1), .I0 (\fsm_output(12)  ), .I1 (nx8012z2), .I2 (
         nx56495z3), .I3 (nx64941z2), .I4 (nx8012z3), .I5 (nx8012z4)) ;
         defparam ix8012z1444.INIT = 64'h0082008200000082;
    LUT5 ix29305z1305 (.O (nx29305z2), .I0 (nx8012z2), .I1 (nx56495z3), .I2 (
         nx64941z2), .I3 (nx8012z3), .I4 (nx8012z4)) ;
         defparam ix29305z1305.INIT = 32'hF6F6FFF6;
    LUT6 ix8012z62810 (.O (nx8012z4), .I0 (p_nbus_image_net_rsc_addr_1_0[13]), .I1 (
         p_nbus_depth_rsc_addr_1_0[2]), .I2 (\fsm_output(12)  ), .I3 (nx56495z5)
         , .I4 (nx1399z2), .I5 (nx56495z4)) ;
         defparam ix8012z62810.INIT = 64'h00F0F0FFC0FAF035;
    (* HLUTNM = "LUT62_1_93" *)
    LUT2 ix9009z1328 (.O (nx9009z1), .I0 (p_image_net_rsc_triosy_lz_1_0), .I1 (
         p_rst_int)) ;
         defparam ix9009z1328.INIT = 4'hE;
    LUT6 ix8049z45004 (.O (nx8049z1), .I0 (nx8049z2), .I1 (nx9046z2), .I2 (
         nx10043z2), .I3 (nx11040z2), .I4 (nx12037z2), .I5 (nx13034z3)) ;
         defparam ix8049z45004.INIT = 64'h6AAAAAAAAAAAAAAA;
    (* HLUTNM = "LUT62_1_28" *)
    LUT5 ix9046z45004 (.O (nx9046z1), .I0 (nx9046z2), .I1 (nx10043z2), .I2 (
         nx11040z2), .I3 (nx12037z2), .I4 (nx13034z3)) ;
         defparam ix9046z45004.INIT = 32'h6AAAAAAA;
    (* HLUTNM = "LUT62_1_28" *)
    LUT4 ix10043z28620 (.O (nx10043z1), .I0 (nx10043z2), .I1 (nx11040z2), .I2 (
         nx12037z2), .I3 (nx13034z3)) ;
         defparam ix10043z28620.INIT = 16'h6AAA;
    (* HLUTNM = "LUT62_1_78" *)
    LUT3 ix11040z1420 (.O (nx11040z1), .I0 (nx11040z2), .I1 (nx12037z2), .I2 (
         nx13034z3)) ;
         defparam ix11040z1420.INIT = 8'h6A;
    (* HLUTNM = "LUT62_1_100" *)
    LUT2 ix12037z1320 (.O (nx12037z1), .I0 (nx12037z2), .I1 (nx13034z3)) ;
         defparam ix12037z1320.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_84" *)
    LUT2 ix40352z1318 (.O (nx40352z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[22])) ;
         defparam ix40352z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_84" *)
    LUT2 ix41349z1318 (.O (nx41349z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[21])) ;
         defparam ix41349z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_83" *)
    LUT2 ix42346z1318 (.O (nx42346z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[20])) ;
         defparam ix42346z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_82" *)
    LUT2 ix43343z1318 (.O (nx43343z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[19])) ;
         defparam ix43343z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_81" *)
    LUT2 ix44340z1319 (.O (nx44340z2), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[18])) ;
         defparam ix44340z1319.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_80" *)
    LUT2 ix45337z1318 (.O (nx45337z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[17])) ;
         defparam ix45337z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_79" *)
    LUT2 ix46334z1318 (.O (nx46334z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[16])) ;
         defparam ix46334z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_74" *)
    LUT2 ix47331z1318 (.O (nx47331z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[15])) ;
         defparam ix47331z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_91" *)
    LUT2 ix48328z1318 (.O (nx48328z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[14])) ;
         defparam ix48328z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_79" *)
    LUT2 ix49325z1318 (.O (nx49325z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[13])) ;
         defparam ix49325z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_93" *)
    LUT2 ix55707z1318 (.O (nx55707z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[12])) ;
         defparam ix55707z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_92" *)
    LUT2 ix54710z1318 (.O (nx54710z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[11])) ;
         defparam ix54710z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_85" *)
    LUT2 ix53713z1318 (.O (nx53713z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[10])) ;
         defparam ix53713z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_83" *)
    LUT2 ix52716z1318 (.O (nx52716z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[9])) ;
         defparam ix52716z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_80" *)
    LUT2 ix51719z1318 (.O (nx51719z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[8])) ;
         defparam ix51719z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_94" *)
    LUT2 ix50722z1318 (.O (nx50722z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[7])) ;
         defparam ix50722z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_81" *)
    LUT2 ix49725z1318 (.O (nx49725z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[6])) ;
         defparam ix49725z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_82" *)
    LUT2 ix48728z1318 (.O (nx48728z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[5])) ;
         defparam ix48728z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_95" *)
    LUT2 ix47731z1318 (.O (nx47731z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[4])) ;
         defparam ix47731z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_96" *)
    LUT2 ix46734z1318 (.O (nx46734z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[3])) ;
         defparam ix46734z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_97" *)
    LUT2 ix44738z1318 (.O (nx44738z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[2])) ;
         defparam ix44738z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_99" *)
    LUT2 ix43741z1318 (.O (nx43741z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[1])) ;
         defparam ix43741z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_101" *)
    LUT2 ix42744z1318 (.O (nx42744z1), .I0 (\fsm_output(6)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0])) ;
         defparam ix42744z1318.INIT = 4'h4;
    (* HLUTNM = "LUT62_1_58" *)
    LUT2 ix44340z1327 (.O (nx44340z1), .I0 (\fsm_output(8)  ), .I1 (
         \fsm_output(6)  )) ;
         defparam ix44340z1327.INIT = 4'hD;
    (* HLUTNM = "LUT62_1_47" *)
    LUT3 ix4577z1523 (.O (nx4577z1), .I0 (p_nbus_depth_rsc_addr_1_0[0]), .I1 (
         \fsm_output(9)  ), .I2 (main_core_inst_z_out_8[8])) ;
         defparam ix4577z1523.INIT = 8'hD1;
    (* HLUTNM = "LUT62_1_47" *)
    LUT4 ix5574z65067 (.O (nx5574z1), .I0 (p_nbus_depth_rsc_addr_1_0[1]), .I1 (
         p_nbus_depth_rsc_addr_1_0[0]), .I2 (\fsm_output(9)  ), .I3 (
         main_core_inst_z_out_8[7])) ;
         defparam ix5574z65067.INIT = 16'hF909;
    LUT5 ix6571z1400 (.O (nx6571z1), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \fsm_output(9)  ), .I4 (main_core_inst_z_out_8[6])) ;
         defparam ix6571z1400.INIT = 32'hFF560056;
    LUT6 ix7568z1482 (.O (nx7568z1), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \fsm_output(9)  ), .I4 (main_core_inst_z_out_8[5]), .I5 (nx1399z3)) ;
         defparam ix7568z1482.INIT = 64'hFF570057FFA800A8;
    LUT6 ix8565z46854 (.O (nx8565z1), .I0 (\fsm_output(9)  ), .I1 (
         \for_1_i_7_0_sva_4(4)  ), .I2 (main_core_inst_z_out_8[4]), .I3 (
         nx1399z3), .I4 (nx7976z4), .I5 (nx7975z4)) ;
         defparam ix8565z46854.INIT = 64'hF5A0F5E4A0A0B1E4;
    LUT6 ix9562z64194 (.O (nx9562z1), .I0 (\fsm_output(9)  ), .I1 (
         \for_1_i_7_0_sva_4(4)  ), .I2 (main_core_inst_z_out_8[3]), .I3 (
         nx64941z4), .I4 (nx1399z3), .I5 (nx7975z4)) ;
         defparam ix9562z64194.INIT = 64'hE4B1F5A0B1E4F5A0;
    LUT6 ix10559z36346 (.O (nx10559z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_z_out_8[2]), .I2 (nx7976z4), .I3 (nx7974z5), .I4 (
         nx7975z8), .I5 (nx7976z5)) ;
         defparam ix10559z36346.INIT = 64'hDDDDDD8D888888D8;
    LUT6 ix11556z36266 (.O (nx11556z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_z_out_8[1]), .I2 (nx7976z4), .I3 (nx7976z5), .I4 (
         nx7977z4), .I5 (nx7977z5)) ;
         defparam ix11556z36266.INIT = 64'hDD8DDDDD88D88888;
    (* HLUTNM = "LUT62_1_63" *)
    LUT2 ix12553z1322 (.O (nx12553z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_z_out_8[0])) ;
         defparam ix12553z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_73" *)
    LUT2 ix13550z1322 (.O (nx13550z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[22])) ;
         defparam ix13550z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_69" *)
    LUT2 ix59274z1322 (.O (nx59274z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[21])) ;
         defparam ix59274z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_61" *)
    LUT2 ix60271z1322 (.O (nx60271z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[20])) ;
         defparam ix60271z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_72" *)
    LUT2 ix61268z1322 (.O (nx61268z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[19])) ;
         defparam ix61268z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_68" *)
    LUT2 ix62265z1322 (.O (nx62265z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[18])) ;
         defparam ix62265z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_64" *)
    LUT2 ix63262z1322 (.O (nx63262z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[17])) ;
         defparam ix63262z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_57" *)
    LUT2 ix64259z1322 (.O (nx64259z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[16])) ;
         defparam ix64259z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_54" *)
    LUT2 ix65256z1322 (.O (nx65256z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[15])) ;
         defparam ix65256z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_60" *)
    LUT2 ix717z1322 (.O (nx717z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[14])) ;
         defparam ix717z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_62" *)
    LUT2 ix1714z1322 (.O (nx1714z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[13])) ;
         defparam ix1714z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_66" *)
    LUT2 ix2711z1322 (.O (nx2711z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[12])) ;
         defparam ix2711z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_65" *)
    LUT2 ix4707z1322 (.O (nx4707z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[11])) ;
         defparam ix4707z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_85" *)
    LUT2 ix5704z1322 (.O (nx5704z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[10])) ;
         defparam ix5704z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_86" *)
    LUT2 ix6701z1322 (.O (nx6701z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[9])) ;
         defparam ix6701z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_101" *)
    LUT2 ix7698z1322 (.O (nx7698z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[8])) ;
         defparam ix7698z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_67" *)
    LUT2 ix8695z1322 (.O (nx8695z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[7])) ;
         defparam ix8695z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_70" *)
    LUT2 ix9692z1322 (.O (nx9692z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[6])) ;
         defparam ix9692z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_71" *)
    LUT2 ix10689z1322 (.O (nx10689z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[5])) ;
         defparam ix10689z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_86" *)
    LUT2 ix11686z1322 (.O (nx11686z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[4])) ;
         defparam ix11686z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_95" *)
    LUT2 ix12683z1322 (.O (nx12683z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[3])) ;
         defparam ix12683z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_96" *)
    LUT2 ix13680z1322 (.O (nx13680z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[2])) ;
         defparam ix13680z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_97" *)
    LUT2 ix15676z1322 (.O (nx15676z1), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[1])) ;
         defparam ix15676z1322.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_102" *)
    LUT2 ix16673z1323 (.O (nx16673z2), .I0 (\fsm_output(9)  ), .I1 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0])) ;
         defparam ix16673z1323.INIT = 4'h8;
    (* HLUTNM = "LUT62_1_59" *)
    LUT2 ix16673z1328 (.O (nx16673z1), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  )) ;
         defparam ix16673z1328.INIT = 4'hE;
    (* HLUTNM = "LUT62_1_74" *)
    LUT4 ix13034z1315 (.O (nx13034z1), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (\fsm_output(6)  ), .I3 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix13034z1315.INIT = 16'h0001;
    (* HLUTNM = "LUT62_1_94" *)
    LUT2 ix63474z1328 (.O (nx63474z1), .I0 (\fsm_output(12)  ), .I1 (
         \fsm_output(4)  )) ;
         defparam ix63474z1328.INIT = 4'hE;
    (* HLUTNM = "LUT62_1_53" *)
    LUT3 ix65061z1316 (.O (nx65061z1), .I0 (nx65061z2), .I1 (\fsm_output(4)  ), 
         .I2 (\fsm_output(0)  )) ;
         defparam ix65061z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_52" *)
    LUT3 ix522z1316 (.O (nx522z1), .I0 (nx522z2), .I1 (\fsm_output(4)  ), .I2 (
         \fsm_output(0)  )) ;
         defparam ix522z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_53" *)
    LUT3 ix1519z1316 (.O (nx1519z1), .I0 (nx1519z2), .I1 (\fsm_output(4)  ), .I2 (
         \fsm_output(0)  )) ;
         defparam ix1519z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_51" *)
    LUT3 ix2516z1316 (.O (nx2516z1), .I0 (nx2516z2), .I1 (\fsm_output(4)  ), .I2 (
         \fsm_output(0)  )) ;
         defparam ix2516z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_91" *)
    LUT3 ix3513z1316 (.O (nx3513z1), .I0 (nx3513z2), .I1 (\fsm_output(4)  ), .I2 (
         \fsm_output(0)  )) ;
         defparam ix3513z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_52" *)
    LUT3 ix4510z1316 (.O (nx4510z1), .I0 (nx4510z2), .I1 (\fsm_output(4)  ), .I2 (
         \fsm_output(0)  )) ;
         defparam ix4510z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_51" *)
    LUT3 ix5507z1316 (.O (nx5507z1), .I0 (nx5507z2), .I1 (\fsm_output(4)  ), .I2 (
         \fsm_output(0)  )) ;
         defparam ix5507z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_50" *)
    LUT3 ix6504z1316 (.O (nx6504z1), .I0 (nx6504z2), .I1 (\fsm_output(4)  ), .I2 (
         \fsm_output(0)  )) ;
         defparam ix6504z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_50" *)
    LUT3 ix7501z1316 (.O (nx7501z1), .I0 (nx7501z2), .I1 (\fsm_output(4)  ), .I2 (
         \fsm_output(0)  )) ;
         defparam ix7501z1316.INIT = 8'h02;
    (* HLUTNM = "LUT62_1_26" *)
    LUT4 ix61860z9557 (.O (nx61860z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[31]), .I3 (
         nx62344z2)) ;
         defparam ix61860z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_23" *)
    LUT4 ix60863z9557 (.O (nx60863z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[30]), .I3 (
         nx63341z2)) ;
         defparam ix60863z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_22" *)
    LUT4 ix59866z9557 (.O (nx59866z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[29]), .I3 (
         nx64338z2)) ;
         defparam ix59866z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_21" *)
    LUT4 ix58869z9557 (.O (nx58869z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[28]), .I3 (
         nx65335z2)) ;
         defparam ix58869z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_20" *)
    LUT4 ix57872z9557 (.O (nx57872z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[27]), .I3 (nx796z2)
         ) ;
         defparam ix57872z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_19" *)
    LUT4 ix56875z9557 (.O (nx56875z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[26]), .I3 (nx1793z2
         )) ;
         defparam ix56875z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_18" *)
    LUT4 ix55878z9557 (.O (nx55878z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[25]), .I3 (nx2790z2
         )) ;
         defparam ix55878z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_17" *)
    LUT4 ix54881z9557 (.O (nx54881z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[24]), .I3 (nx3787z2
         )) ;
         defparam ix54881z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_15" *)
    LUT4 ix53884z9557 (.O (nx53884z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[23]), .I3 (nx4784z2
         )) ;
         defparam ix53884z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_14" *)
    LUT4 ix52887z9557 (.O (nx52887z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[22]), .I3 (nx5781z2
         )) ;
         defparam ix52887z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_13" *)
    LUT4 ix52591z9557 (.O (nx52591z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[21]), .I3 (
         nx46829z2)) ;
         defparam ix52591z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_12" *)
    LUT4 ix51594z9557 (.O (nx51594z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[20]), .I3 (
         nx47826z2)) ;
         defparam ix51594z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_11" *)
    LUT4 ix50597z9557 (.O (nx50597z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[19]), .I3 (
         nx48823z2)) ;
         defparam ix50597z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_10" *)
    LUT4 ix49600z9557 (.O (nx49600z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[18]), .I3 (
         nx49820z2)) ;
         defparam ix49600z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_9" *)
    LUT4 ix48603z9557 (.O (nx48603z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[17]), .I3 (
         nx50817z2)) ;
         defparam ix48603z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_8" *)
    LUT4 ix47606z9557 (.O (nx47606z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[16]), .I3 (
         nx51814z2)) ;
         defparam ix47606z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_7" *)
    LUT4 ix46609z9557 (.O (nx46609z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[15]), .I3 (
         nx52811z2)) ;
         defparam ix46609z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_5" *)
    LUT4 ix45612z9557 (.O (nx45612z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[14]), .I3 (
         nx53808z2)) ;
         defparam ix45612z9557.INIT = 16'h2033;
    LUT4 ix44615z9557 (.O (nx44615z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[13]), .I3 (
         nx54805z2)) ;
         defparam ix44615z9557.INIT = 16'h2033;
    LUT4 ix43618z9557 (.O (nx43618z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[12]), .I3 (
         nx55802z2)) ;
         defparam ix43618z9557.INIT = 16'h2033;
    LUT4 ix41622z9557 (.O (nx41622z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[11]), .I3 (
         nx57798z2)) ;
         defparam ix41622z9557.INIT = 16'h2033;
    LUT4 ix40625z9557 (.O (nx40625z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[10]), .I3 (
         nx58795z2)) ;
         defparam ix40625z9557.INIT = 16'h2033;
    LUT4 ix39628z9557 (.O (nx39628z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[9]), .I3 (nx59792z2
         )) ;
         defparam ix39628z9557.INIT = 16'h2033;
    LUT4 ix38631z9557 (.O (nx38631z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[8]), .I3 (nx60789z2
         )) ;
         defparam ix38631z9557.INIT = 16'h2033;
    LUT4 ix37634z9557 (.O (nx37634z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[7]), .I3 (nx61786z2
         )) ;
         defparam ix37634z9557.INIT = 16'h2033;
    LUT4 ix36637z9557 (.O (nx36637z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[6]), .I3 (nx62783z2
         )) ;
         defparam ix36637z9557.INIT = 16'h2033;
    LUT4 ix35640z9557 (.O (nx35640z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[5]), .I3 (nx63780z2
         )) ;
         defparam ix35640z9557.INIT = 16'h2033;
    LUT4 ix34643z9557 (.O (nx34643z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[4]), .I3 (nx64777z2
         )) ;
         defparam ix34643z9557.INIT = 16'h2033;
    LUT4 ix33646z9557 (.O (nx33646z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[3]), .I3 (nx238z2)
         ) ;
         defparam ix33646z9557.INIT = 16'h2033;
    LUT4 ix32649z9557 (.O (nx32649z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[2]), .I3 (nx1235z2)
         ) ;
         defparam ix32649z9557.INIT = 16'h2033;
    LUT4 ix30653z9557 (.O (nx30653z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[1]), .I3 (nx3231z2)
         ) ;
         defparam ix30653z9557.INIT = 16'h2033;
    LUT4 ix29656z9557 (.O (nx29656z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[0]), .I3 (nx4228z2)
         ) ;
         defparam ix29656z9557.INIT = 16'h2033;
    (* HLUTNM = "LUT62_1_26" *)
    LUT5 ix62344z14421 (.O (nx62344z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[31]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx62344z2)) ;
         defparam ix62344z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_58" *)
    LUT4 ix62344z6274 (.O (nx62344z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[31]), .I3 (
         main_core_inst_z_out_6[0])) ;
         defparam ix62344z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_23" *)
    LUT5 ix63341z14421 (.O (nx63341z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[30]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx63341z2)) ;
         defparam ix63341z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_59" *)
    LUT4 ix63341z6274 (.O (nx63341z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[30]), .I3 (
         main_core_inst_z_out_6[1])) ;
         defparam ix63341z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_22" *)
    LUT5 ix64338z14421 (.O (nx64338z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[29]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx64338z2)) ;
         defparam ix64338z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_60" *)
    LUT4 ix64338z6274 (.O (nx64338z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[29]), .I3 (
         main_core_inst_z_out_6[2])) ;
         defparam ix64338z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_21" *)
    LUT5 ix65335z14421 (.O (nx65335z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[28]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx65335z2)) ;
         defparam ix65335z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_54" *)
    LUT4 ix65335z6274 (.O (nx65335z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[28]), .I3 (
         main_core_inst_z_out_6[3])) ;
         defparam ix65335z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_20" *)
    LUT5 ix796z14421 (.O (nx796z1), .I0 (\fsm_output(6)  ), .I1 (\fsm_output(5)  
         ), .I2 (main_core_inst_reconstruction_error_rec_error_lpi_6[27]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx796z2)) ;
         defparam ix796z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_61" *)
    LUT4 ix796z6274 (.O (nx796z2), .I0 (\fsm_output(9)  ), .I1 (\fsm_output(8)  
         ), .I2 (main_core_inst_reconstruction_error_rec_error_sva[27]), .I3 (
         main_core_inst_z_out_6[4])) ;
         defparam ix796z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_19" *)
    LUT5 ix1793z14421 (.O (nx1793z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[26]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx1793z2)) ;
         defparam ix1793z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_62" *)
    LUT4 ix1793z6274 (.O (nx1793z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[26]), .I3 (
         main_core_inst_z_out_6[5])) ;
         defparam ix1793z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_18" *)
    LUT5 ix2790z14421 (.O (nx2790z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[25]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx2790z2)) ;
         defparam ix2790z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_63" *)
    LUT4 ix2790z6274 (.O (nx2790z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[25]), .I3 (
         main_core_inst_z_out_6[6])) ;
         defparam ix2790z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_17" *)
    LUT5 ix3787z14421 (.O (nx3787z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[24]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx3787z2)) ;
         defparam ix3787z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_64" *)
    LUT4 ix3787z6274 (.O (nx3787z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[24]), .I3 (
         main_core_inst_z_out_6[7])) ;
         defparam ix3787z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_15" *)
    LUT5 ix4784z14421 (.O (nx4784z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[23]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx4784z2)) ;
         defparam ix4784z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_65" *)
    LUT4 ix4784z6274 (.O (nx4784z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[23]), .I3 (
         main_core_inst_z_out_6[8])) ;
         defparam ix4784z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_14" *)
    LUT5 ix5781z14421 (.O (nx5781z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[22]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx5781z2)) ;
         defparam ix5781z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_66" *)
    LUT4 ix5781z6274 (.O (nx5781z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[22]), .I3 (
         main_core_inst_z_out_6[9])) ;
         defparam ix5781z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_13" *)
    LUT5 ix46829z14421 (.O (nx46829z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[21]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx46829z2)) ;
         defparam ix46829z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_67" *)
    LUT4 ix46829z6274 (.O (nx46829z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[21]), .I3 (
         main_core_inst_z_out_6[10])) ;
         defparam ix46829z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_12" *)
    LUT5 ix47826z14421 (.O (nx47826z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[20]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx47826z2)) ;
         defparam ix47826z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_68" *)
    LUT4 ix47826z6274 (.O (nx47826z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[20]), .I3 (
         main_core_inst_z_out_6[11])) ;
         defparam ix47826z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_11" *)
    LUT5 ix48823z14421 (.O (nx48823z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[19]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx48823z2)) ;
         defparam ix48823z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_69" *)
    LUT4 ix48823z6274 (.O (nx48823z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[19]), .I3 (
         main_core_inst_z_out_6[12])) ;
         defparam ix48823z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_10" *)
    LUT5 ix49820z14421 (.O (nx49820z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[18]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx49820z2)) ;
         defparam ix49820z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_70" *)
    LUT4 ix49820z6274 (.O (nx49820z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[18]), .I3 (
         main_core_inst_z_out_6[13])) ;
         defparam ix49820z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_9" *)
    LUT5 ix50817z14421 (.O (nx50817z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[17]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx50817z2)) ;
         defparam ix50817z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_71" *)
    LUT4 ix50817z6274 (.O (nx50817z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[17]), .I3 (
         main_core_inst_z_out_6[14])) ;
         defparam ix50817z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_8" *)
    LUT5 ix51814z14421 (.O (nx51814z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[16]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx51814z2)) ;
         defparam ix51814z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_72" *)
    LUT4 ix51814z6274 (.O (nx51814z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[16]), .I3 (
         main_core_inst_z_out_6[15])) ;
         defparam ix51814z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_7" *)
    LUT5 ix52811z14421 (.O (nx52811z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[15]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx52811z2)) ;
         defparam ix52811z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_73" *)
    LUT4 ix52811z6274 (.O (nx52811z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[15]), .I3 (
         main_core_inst_z_out_6[16])) ;
         defparam ix52811z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_5" *)
    LUT5 ix53808z14421 (.O (nx53808z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[14]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx53808z2)) ;
         defparam ix53808z14421.INIT = 32'h30203333;
    (* HLUTNM = "LUT62_1_57" *)
    LUT4 ix53808z6274 (.O (nx53808z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[14]), .I3 (
         main_core_inst_z_out_6[17])) ;
         defparam ix53808z6274.INIT = 16'h135F;
    LUT5 ix54805z14421 (.O (nx54805z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[13]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx54805z2)) ;
         defparam ix54805z14421.INIT = 32'h30203333;
    LUT4 ix54805z6274 (.O (nx54805z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[13]), .I3 (
         main_core_inst_z_out_6[18])) ;
         defparam ix54805z6274.INIT = 16'h135F;
    LUT5 ix55802z14421 (.O (nx55802z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[12]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx55802z2)) ;
         defparam ix55802z14421.INIT = 32'h30203333;
    LUT4 ix55802z6274 (.O (nx55802z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[12]), .I3 (
         main_core_inst_z_out_6[19])) ;
         defparam ix55802z6274.INIT = 16'h135F;
    LUT5 ix57798z14421 (.O (nx57798z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[11]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx57798z2)) ;
         defparam ix57798z14421.INIT = 32'h30203333;
    LUT4 ix57798z6274 (.O (nx57798z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[11]), .I3 (
         main_core_inst_z_out_6[20])) ;
         defparam ix57798z6274.INIT = 16'h135F;
    LUT5 ix58795z14421 (.O (nx58795z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[10]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx58795z2)) ;
         defparam ix58795z14421.INIT = 32'h30203333;
    LUT4 ix58795z6274 (.O (nx58795z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[10]), .I3 (
         main_core_inst_z_out_6[21])) ;
         defparam ix58795z6274.INIT = 16'h135F;
    LUT5 ix59792z14421 (.O (nx59792z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[9]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx59792z2)) ;
         defparam ix59792z14421.INIT = 32'h30203333;
    LUT4 ix59792z6274 (.O (nx59792z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[9]), .I3 (
         main_core_inst_z_out_6[22])) ;
         defparam ix59792z6274.INIT = 16'h135F;
    LUT5 ix60789z14421 (.O (nx60789z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[8]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx60789z2)) ;
         defparam ix60789z14421.INIT = 32'h30203333;
    LUT4 ix60789z6274 (.O (nx60789z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[8]), .I3 (
         main_core_inst_z_out_6[23])) ;
         defparam ix60789z6274.INIT = 16'h135F;
    LUT5 ix61786z14421 (.O (nx61786z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[7]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx61786z2)) ;
         defparam ix61786z14421.INIT = 32'h30203333;
    LUT4 ix61786z6274 (.O (nx61786z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[7]), .I3 (
         main_core_inst_z_out_6[24])) ;
         defparam ix61786z6274.INIT = 16'h135F;
    LUT5 ix62783z14421 (.O (nx62783z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[6]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx62783z2)) ;
         defparam ix62783z14421.INIT = 32'h30203333;
    LUT4 ix62783z6274 (.O (nx62783z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[6]), .I3 (
         main_core_inst_z_out_6[25])) ;
         defparam ix62783z6274.INIT = 16'h135F;
    LUT5 ix63780z14421 (.O (nx63780z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[5]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx63780z2)) ;
         defparam ix63780z14421.INIT = 32'h30203333;
    LUT4 ix63780z6274 (.O (nx63780z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[5]), .I3 (
         main_core_inst_z_out_6[26])) ;
         defparam ix63780z6274.INIT = 16'h135F;
    LUT5 ix64777z14421 (.O (nx64777z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[4]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx64777z2)) ;
         defparam ix64777z14421.INIT = 32'h30203333;
    LUT4 ix64777z6274 (.O (nx64777z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[4]), .I3 (
         main_core_inst_z_out_6[27])) ;
         defparam ix64777z6274.INIT = 16'h135F;
    LUT5 ix238z14421 (.O (nx238z1), .I0 (\fsm_output(6)  ), .I1 (\fsm_output(5)  
         ), .I2 (main_core_inst_reconstruction_error_rec_error_lpi_6[3]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx238z2)) ;
         defparam ix238z14421.INIT = 32'h30203333;
    LUT4 ix238z6274 (.O (nx238z2), .I0 (\fsm_output(9)  ), .I1 (\fsm_output(8)  
         ), .I2 (main_core_inst_reconstruction_error_rec_error_sva[3]), .I3 (
         main_core_inst_z_out_6[28])) ;
         defparam ix238z6274.INIT = 16'h135F;
    LUT5 ix1235z14421 (.O (nx1235z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[2]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx1235z2)) ;
         defparam ix1235z14421.INIT = 32'h30203333;
    LUT4 ix1235z6274 (.O (nx1235z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[2]), .I3 (
         main_core_inst_z_out_6[29])) ;
         defparam ix1235z6274.INIT = 16'h135F;
    LUT5 ix3231z14421 (.O (nx3231z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[1]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx3231z2)) ;
         defparam ix3231z14421.INIT = 32'h30203333;
    LUT4 ix3231z6274 (.O (nx3231z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[1]), .I3 (
         main_core_inst_z_out_6[30])) ;
         defparam ix3231z6274.INIT = 16'h135F;
    LUT5 ix4228z14421 (.O (nx4228z1), .I0 (\fsm_output(6)  ), .I1 (
         \fsm_output(5)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[0]), .I3 (
         \p_for_for_mux1h_2_nl(1)  ), .I4 (nx4228z2)) ;
         defparam ix4228z14421.INIT = 32'h30203333;
    LUT4 ix4228z6274 (.O (nx4228z2), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(8)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I3 (
         main_core_inst_z_out_6[31])) ;
         defparam ix4228z6274.INIT = 16'h135F;
    (* HLUTNM = "LUT62_1_46" *)
    LUT3 ix56642z1341 (.O (nx56642z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[8]), .I2 (nx56642z2)) ;
         defparam ix56642z1341.INIT = 8'h1B;
    (* HLUTNM = "LUT62_1_16" *)
    LUT5 ix57639z49974 (.O (nx57639z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[8]), .I3 (nx57639z2), .I4 (nx56642z2
         )) ;
         defparam ix57639z49974.INIT = 32'h14BEBE14;
    LUT6 ix27832z62310 (.O (nx27832z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[0]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[8]), .I3 (nx11510z4), .I4 (nx56642z2
         ), .I5 (nx27832z2)) ;
         defparam ix27832z62310.INIT = 64'h14BEBE14EE44EE44;
    (* HLUTNM = "LUT62_1_16" *)
    LUT4 ix11510z59685 (.O (nx11510z6), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I2 (nx57639z2), .I3 (nx56642z2
         )) ;
         defparam ix11510z59685.INIT = 16'hE400;
    (* HLUTNM = "LUT62_1_39" *)
    LUT4 ix11510z6504 (.O (nx11510z5), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[0]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I3 (
         main_core_inst_for_for_j_8_0_sva_3[8])) ;
         defparam ix11510z6504.INIT = 16'h1444;
    LUT6 ix26835z62310 (.O (nx26835z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[1]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[8]), .I3 (nx13034z3), .I4 (nx56642z2
         ), .I5 (nx26835z2)) ;
         defparam ix26835z62310.INIT = 64'h14BEBE14EE44EE44;
    (* HLUTNM = "LUT62_1_32" *)
    LUT5 ix26835z17763 (.O (nx26835z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[0]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I3 (nx11510z4), .I4 (nx57639z2
         )) ;
         defparam ix26835z17763.INIT = 32'hEA404040;
    LUT6 ix25838z59910 (.O (nx25838z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[2]), .I2 (nx12037z2), .I3 (nx25838z2
         ), .I4 (nx25838z3), .I5 (nx25838z4)) ;
         defparam ix25838z59910.INIT = 64'hE41BE4E4E4E4E4E4;
    LUT6 ix24841z1313 (.O (nx24841z1), .I0 (nx25838z2), .I1 (nx25838z3), .I2 (
         nx25838z4), .I3 (nx24841z2), .I4 (nx24841z3), .I5 (nx24841z4)) ;
         defparam ix24841z1313.INIT = 64'h0000BFFF4000FFFF;
    (* HLUTNM = "LUT62_1_76" *)
    LUT3 ix24841z1545 (.O (nx24841z4), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (nx11040z2)) ;
         defparam ix24841z1545.INIT = 8'hE4;
    (* HLUTNM = "LUT62_1_31" *)
    LUT3 ix24841z1343 (.O (nx24841z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (nx11040z2)) ;
         defparam ix24841z1343.INIT = 8'h1B;
    (* HLUTNM = "LUT62_1_78" *)
    LUT3 ix24841z1543 (.O (nx24841z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[2]), .I2 (nx12037z2)) ;
         defparam ix24841z1543.INIT = 8'hE4;
    LUT4 ix23844z8454 (.O (nx23844z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I2 (nx10043z2), .I3 (nx23844z2
         )) ;
         defparam ix23844z8454.INIT = 16'h1BE4;
    (* HLUTNM = "LUT62_1_25" *)
    LUT5 ix11514z23161 (.O (nx11514z4), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I1 (nx25838z2), .I2 (nx25838z3
         ), .I3 (nx25838z4), .I4 (nx23844z3)) ;
         defparam ix11514z23161.INIT = 32'h65555555;
    LUT6 ix11514z36267 (.O (nx11514z3), .I0 (\p_fsm_output(10)  ), .I1 (
         nx10043z2), .I2 (nx25838z2), .I3 (nx25838z3), .I4 (nx25838z4), .I5 (
         nx23844z3)) ;
         defparam ix11514z36267.INIT = 64'h8288888888888888;
    LUT6 ix22847z62310 (.O (nx22847z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I3 (nx9046z2), .I4 (nx10043z2)
         , .I5 (nx23844z2)) ;
         defparam ix22847z62310.INIT = 64'h14BEBE14EE44EE44;
    LUT6 ix11515z23161 (.O (nx11515z4), .I0 (nx9046z2), .I1 (nx10043z2), .I2 (
         nx25838z2), .I3 (nx25838z3), .I4 (nx25838z4), .I5 (nx23844z3)) ;
         defparam ix11515z23161.INIT = 64'h5955555555555555;
    LUT6 ix11515z23160 (.O (nx11515z3), .I0 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I2 (nx25838z2), .I3 (nx25838z3
         ), .I4 (nx25838z4), .I5 (nx23844z3)) ;
         defparam ix11515z23160.INIT = 64'h5955555555555555;
    LUT6 ix21850z1569 (.O (nx21850z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I3 (nx21850z2), .I4 (nx23844z2
         ), .I5 (nx21850z3)) ;
         defparam ix21850z1569.INIT = 64'hEA1500FF00FF00FF;
    LUT6 ix11516z1318 (.O (nx11516z6), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[6]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I3 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I4 (nx8049z2), .I5 (nx21850z3)
         ) ;
         defparam ix11516z1318.INIT = 64'h1000BAAA00000000;
    LUT6 ix11516z23161 (.O (nx11516z4), .I0 (nx21850z2), .I1 (nx25838z2), .I2 (
         nx25838z3), .I3 (nx25838z4), .I4 (nx23844z3), .I5 (nx11516z5)) ;
         defparam ix11516z23161.INIT = 64'h4555555555555555;
    (* HLUTNM = "LUT62_1_2" *)
    LUT5 ix11516z17765 (.O (nx11516z5), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I3 (nx9046z2), .I4 (nx10043z2)
         ) ;
         defparam ix11516z17765.INIT = 32'hEA404040;
    (* HLUTNM = "LUT62_1_2" *)
    LUT5 ix21850z17764 (.O (nx21850z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I3 (nx9046z2), .I4 (nx10043z2)
         ) ;
         defparam ix21850z17764.INIT = 32'hFF404040;
    (* HLUTNM = "LUT62_1_25" *)
    LUT4 ix23844z3363 (.O (nx23844z2), .I0 (nx23844z3), .I1 (nx25838z4), .I2 (
         nx25838z2), .I3 (nx25838z3)) ;
         defparam ix23844z3363.INIT = 16'h0800;
    (* HLUTNM = "LUT62_1_31" *)
    LUT5 ix23844z17764 (.O (nx23844z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[2]), .I3 (nx11040z2), .I4 (nx12037z2
         )) ;
         defparam ix23844z17764.INIT = 32'hEA404040;
    LUT5 ix25838z17765 (.O (nx25838z4), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[1]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[0]), .I3 (nx13034z3), .I4 (nx11510z4
         )) ;
         defparam ix25838z17765.INIT = 32'hFF404040;
    (* HLUTNM = "LUT62_1_46" *)
    LUT4 ix25838z59752 (.O (nx25838z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I2 (nx57639z2), .I3 (nx56642z2
         )) ;
         defparam ix25838z59752.INIT = 16'hE444;
    (* HLUTNM = "LUT62_1_39" *)
    LUT4 ix25838z6776 (.O (nx25838z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[1]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[0]), .I3 (
         main_core_inst_for_for_j_8_0_sva_3[8])) ;
         defparam ix25838z6776.INIT = 16'h1555;
    (* HLUTNM = "LUT62_1_32" *)
    LUT3 ix27832z1543 (.O (nx27832z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I2 (nx57639z2)) ;
         defparam ix27832z1543.INIT = 8'hE4;
    (* HLUTNM = "LUT62_1_76" *)
    LUT3 ix21850z1342 (.O (nx21850z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[6]), .I2 (nx8049z2)) ;
         defparam ix21850z1342.INIT = 8'h1B;
    (* HLUTNM = "LUT62_1_45" *)
    LUT4 ix5387z14882 (.O (nx5387z1), .I0 (p_nbus_image_net_rsc_addr_1_0[15]), .I1 (
         p_nbus_depth_rsc_addr_1_0[0]), .I2 (\fsm_output(12)  ), .I3 (
         \fsm_output(4)  )) ;
         defparam ix5387z14882.INIT = 16'h3500;
    (* HLUTNM = "LUT62_1_56" *)
    LUT2 ix63474z1319 (.O (nx63474z2), .I0 (p_nbus_depth_rsc_addr_1_0[0]), .I1 (
         \fsm_output(12)  )) ;
         defparam ix63474z1319.INIT = 4'h4;
    LUT6 ix4390z1314 (.O (nx4390z1), .I0 (p_nbus_image_net_rsc_addr_1_0[14]), .I1 (
         p_nbus_image_net_rsc_addr_1_0[15]), .I2 (p_nbus_depth_rsc_addr_1_0[1])
         , .I3 (p_nbus_depth_rsc_addr_1_0[0]), .I4 (\fsm_output(12)  ), .I5 (
         \fsm_output(4)  )) ;
         defparam ix4390z1314.INIT = 64'h0FF0666600000000;
    (* HLUTNM = "LUT62_1_36" *)
    LUT3 ix62477z1354 (.O (nx62477z1), .I0 (\fsm_output(12)  ), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0])) ;
         defparam ix62477z1354.INIT = 8'h28;
    (* HLUTNM = "LUT62_1_33" *)
    LUT5 ix3393z14882 (.O (nx3393z1), .I0 (p_nbus_image_net_rsc_addr_1_0[13]), .I1 (
         p_nbus_depth_rsc_addr_1_0[2]), .I2 (\fsm_output(12)  ), .I3 (
         \fsm_output(4)  ), .I4 (nx56495z4)) ;
         defparam ix3393z14882.INIT = 32'hCA003500;
    LUT6 ix2396z14882 (.O (nx2396z1), .I0 (p_nbus_image_net_rsc_addr_1_0[13]), .I1 (
         p_nbus_depth_rsc_addr_1_0[2]), .I2 (\fsm_output(12)  ), .I3 (
         \fsm_output(4)  ), .I4 (nx1399z2), .I5 (nx56495z4)) ;
         defparam ix2396z14882.INIT = 64'h0000FF00CA003500;
    LUT5 ix1399z10058 (.O (nx1399z1), .I0 (\fsm_output(4)  ), .I1 (nx56495z5), .I2 (
         nx1399z2), .I3 (nx1399z4), .I4 (nx56495z4)) ;
         defparam ix1399z10058.INIT = 32'h22222228;
    LUT6 ix402z10058 (.O (nx402z1), .I0 (\fsm_output(4)  ), .I1 (nx64941z3), .I2 (
         nx56495z5), .I3 (nx1399z2), .I4 (nx1399z4), .I5 (nx56495z4)) ;
         defparam ix402z10058.INIT = 64'h2222222222222228;
    LUT5 ix8012z45005 (.O (nx8012z3), .I0 (nx64941z3), .I1 (nx56495z5), .I2 (
         nx1399z2), .I3 (nx1399z4), .I4 (nx56495z4)) ;
         defparam ix8012z45005.INIT = 32'hAAAAAAA9;
    (* HLUTNM = "LUT62_1_35" *)
    LUT5 ix58489z17763 (.O (nx58489z2), .I0 (\fsm_output(12)  ), .I1 (
         \for_i_7_0_sva_3(4)  ), .I2 (\for_i_7_0_sva_3(3)  ), .I3 (
         \for_1_i_7_0_sva_4(4)  ), .I4 (nx1399z3)) ;
         defparam ix58489z17763.INIT = 32'hEA404040;
    (* HLUTNM = "LUT62_1_98" *)
    LUT2 ix64941z1316 (.O (nx64941z1), .I0 (\fsm_output(4)  ), .I1 (nx64941z2)
         ) ;
         defparam ix64941z1316.INIT = 4'h2;
    LUT6 ix64941z45004 (.O (nx64941z2), .I0 (nx56495z6), .I1 (nx64941z3), .I2 (
         nx56495z5), .I3 (nx1399z2), .I4 (nx1399z4), .I5 (nx56495z4)) ;
         defparam ix64941z45004.INIT = 64'hAAAAAAAAAAAAAAA9;
    (* HLUTNM = "LUT62_1_37" *)
    LUT5 ix63944z52579 (.O (nx63944z2), .I0 (\fsm_output(12)  ), .I1 (
         \fsm_output(4)  ), .I2 (\for_i_7_0_sva_3(7)  ), .I3 (nx63944z3), .I4 (
         nx56495z3)) ;
         defparam ix63944z52579.INIT = 32'h048CC840;
    LUT6 ix56495z1317 (.O (nx56495z3), .I0 (nx56495z4), .I1 (nx56495z5), .I2 (
         nx1399z2), .I3 (nx1399z4), .I4 (nx56495z6), .I5 (nx64941z3)) ;
         defparam ix56495z1317.INIT = 64'h0000000000000001;
    (* HLUTNM = "LUT62_1_36" *)
    LUT5 ix56495z31900 (.O (nx56495z4), .I0 (p_nbus_image_net_rsc_addr_1_0[14])
         , .I1 (p_nbus_image_net_rsc_addr_1_0[15]), .I2 (
         p_nbus_depth_rsc_addr_1_0[1]), .I3 (p_nbus_depth_rsc_addr_1_0[0]), .I4 (
         \fsm_output(12)  )) ;
         defparam ix56495z31900.INIT = 32'h0FFF7777;
    (* HLUTNM = "LUT62_1_33" *)
    LUT3 ix1399z1369 (.O (nx1399z4), .I0 (p_nbus_image_net_rsc_addr_1_0[13]), .I1 (
         p_nbus_depth_rsc_addr_1_0[2]), .I2 (\fsm_output(12)  )) ;
         defparam ix1399z1369.INIT = 8'h35;
    (* HLUTNM = "LUT62_1_75" *)
    LUT3 ix1399z1342 (.O (nx1399z2), .I0 (\fsm_output(12)  ), .I1 (
         \for_i_7_0_sva_3(3)  ), .I2 (nx1399z3)) ;
         defparam ix1399z1342.INIT = 8'h1B;
    (* HLUTNM = "LUT62_1_35" *)
    LUT3 ix56495z1345 (.O (nx56495z5), .I0 (\fsm_output(12)  ), .I1 (
         \for_i_7_0_sva_3(4)  ), .I2 (\for_1_i_7_0_sva_4(4)  )) ;
         defparam ix56495z1345.INIT = 8'h1B;
    (* HLUTNM = "LUT62_1_75" *)
    LUT3 ix64941z1343 (.O (nx64941z3), .I0 (\fsm_output(12)  ), .I1 (
         \for_i_7_0_sva_3(5)  ), .I2 (nx64941z4)) ;
         defparam ix64941z1343.INIT = 8'h1B;
    (* HLUTNM = "LUT62_1_92" *)
    LUT3 ix56495z1346 (.O (nx56495z6), .I0 (\fsm_output(12)  ), .I1 (
         \for_i_7_0_sva_3(6)  ), .I2 (nx56495z7)) ;
         defparam ix56495z1346.INIT = 8'h1B;
    (* HLUTNM = "LUT62_1_37" *)
    LUT3 ix8012z1342 (.O (nx8012z2), .I0 (\fsm_output(12)  ), .I1 (
         \for_i_7_0_sva_3(7)  ), .I2 (nx63944z3)) ;
         defparam ix8012z1342.INIT = 8'h1B;
    (* HLUTNM = "LUT62_1_42" *)
    LUT2 ix63944z1328 (.O (nx63944z1), .I0 (\fsm_output(4)  ), .I1 (
         \fsm_output(0)  )) ;
         defparam ix63944z1328.INIT = 4'hE;
    LUT2 ix42790z1336 (.O (nx42790z15), .I0 (
         p_nbus_image_error_rsc_data_out_int[0]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1336.INIT = 4'h8;
    LUT2 ix42790z1335 (.O (nx42790z14), .I0 (
         p_nbus_image_error_rsc_data_out_int[1]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1335.INIT = 4'h8;
    LUT2 ix42790z1334 (.O (nx42790z13), .I0 (
         p_nbus_image_error_rsc_data_out_int[2]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1334.INIT = 4'h8;
    LUT2 ix42790z1333 (.O (nx42790z12), .I0 (
         p_nbus_image_error_rsc_data_out_int[3]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1333.INIT = 4'h8;
    LUT2 ix42790z1332 (.O (nx42790z11), .I0 (
         p_nbus_image_error_rsc_data_out_int[4]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1332.INIT = 4'h8;
    LUT2 ix42790z1331 (.O (nx42790z10), .I0 (
         p_nbus_image_error_rsc_data_out_int[5]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1331.INIT = 4'h8;
    LUT2 ix42790z1330 (.O (nx42790z9), .I0 (
         p_nbus_image_error_rsc_data_out_int[6]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1330.INIT = 4'h8;
    LUT2 ix42790z1329 (.O (nx42790z8), .I0 (
         p_nbus_image_error_rsc_data_out_int[7]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1329.INIT = 4'h8;
    LUT2 ix42790z1328 (.O (nx42790z7), .I0 (
         p_nbus_image_error_rsc_data_out_int[8]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1328.INIT = 4'h8;
    LUT2 ix42790z1327 (.O (nx42790z6), .I0 (
         p_nbus_image_error_rsc_data_out_int[9]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1327.INIT = 4'h8;
    LUT2 ix42790z1326 (.O (nx42790z5), .I0 (
         p_nbus_image_error_rsc_data_out_int[10]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1326.INIT = 4'h8;
    LUT2 ix42790z1325 (.O (nx42790z4), .I0 (
         p_nbus_image_error_rsc_data_out_int[11]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1325.INIT = 4'h8;
    LUT2 ix42790z1324 (.O (nx42790z3), .I0 (
         p_nbus_image_error_rsc_data_out_int[12]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1324.INIT = 4'h8;
    LUT2 ix42790z1323 (.O (nx42790z2), .I0 (
         p_nbus_image_error_rsc_data_out_int[13]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1323.INIT = 4'h8;
    LUT2 ix42790z1322 (.O (nx42790z1), .I0 (
         p_nbus_image_error_rsc_data_out_int[14]), .I1 (\fsm_output(8)  )) ;
         defparam ix42790z1322.INIT = 4'h8;
    LUT4 ix6176z1330 (.O (nx6176z15), .I0 (
         p_nbus_image_error_rsc_data_out_int[0]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1330.INIT = 16'h0002;
    LUT4 ix6176z1329 (.O (nx6176z14), .I0 (
         p_nbus_image_error_rsc_data_out_int[1]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1329.INIT = 16'h0002;
    LUT4 ix6176z1328 (.O (nx6176z13), .I0 (
         p_nbus_image_error_rsc_data_out_int[2]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1328.INIT = 16'h0002;
    LUT4 ix6176z1327 (.O (nx6176z12), .I0 (
         p_nbus_image_error_rsc_data_out_int[3]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1327.INIT = 16'h0002;
    LUT4 ix6176z1326 (.O (nx6176z11), .I0 (
         p_nbus_image_error_rsc_data_out_int[4]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1326.INIT = 16'h0002;
    LUT4 ix6176z1325 (.O (nx6176z10), .I0 (
         p_nbus_image_error_rsc_data_out_int[5]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1325.INIT = 16'h0002;
    LUT4 ix6176z1324 (.O (nx6176z9), .I0 (p_nbus_image_error_rsc_data_out_int[6]
         ), .I1 (\p_fsm_output(10)  ), .I2 (\fsm_output(1)  ), .I3 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1324.INIT = 16'h0002;
    LUT4 ix6176z1323 (.O (nx6176z8), .I0 (p_nbus_image_error_rsc_data_out_int[7]
         ), .I1 (\p_fsm_output(10)  ), .I2 (\fsm_output(1)  ), .I3 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1323.INIT = 16'h0002;
    LUT4 ix6176z1322 (.O (nx6176z7), .I0 (p_nbus_image_error_rsc_data_out_int[8]
         ), .I1 (\p_fsm_output(10)  ), .I2 (\fsm_output(1)  ), .I3 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1322.INIT = 16'h0002;
    LUT4 ix6176z1321 (.O (nx6176z6), .I0 (p_nbus_image_error_rsc_data_out_int[9]
         ), .I1 (\p_fsm_output(10)  ), .I2 (\fsm_output(1)  ), .I3 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1321.INIT = 16'h0002;
    LUT4 ix6176z1320 (.O (nx6176z5), .I0 (
         p_nbus_image_error_rsc_data_out_int[10]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1320.INIT = 16'h0002;
    LUT4 ix6176z1319 (.O (nx6176z4), .I0 (
         p_nbus_image_error_rsc_data_out_int[11]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1319.INIT = 16'h0002;
    LUT4 ix6176z1318 (.O (nx6176z3), .I0 (
         p_nbus_image_error_rsc_data_out_int[12]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1318.INIT = 16'h0002;
    LUT4 ix6176z1317 (.O (nx6176z2), .I0 (
         p_nbus_image_error_rsc_data_out_int[13]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1317.INIT = 16'h0002;
    LUT4 ix6176z1316 (.O (nx6176z1), .I0 (
         p_nbus_image_error_rsc_data_out_int[14]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix6176z1316.INIT = 16'h0002;
    LUT5 ix10394z1338 (.O (nx10394z43), .I0 (
         p_nbus_image_error_rsc_data_out_int[15]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (\fsm_output(1)  ), .I4 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix10394z1338.INIT = 32'hFFFFFFEC;
    LUT4 ix10394z1393 (.O (nx10394z42), .I0 (
         p_nbus_image_error_rsc_data_out_int[16]), .I1 (\fsm_output(8)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix10394z1393.INIT = 16'hFFF8;
    LUT5 ix10394z1375 (.O (nx10394z40), .I0 (
         p_nbus_image_error_rsc_data_out_int[17]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (\fsm_output(1)  ), .I4 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix10394z1375.INIT = 32'hFFFFFFEC;
    LUT5 ix10394z1332 (.O (nx10394z39), .I0 (
         p_nbus_image_error_rsc_data_out_int[18]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (\fsm_output(1)  ), .I4 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix10394z1332.INIT = 32'hFFFFFFEC;
    LUT2 ix10394z1350 (.O (nx10394z29), .I0 (
         p_nbus_image_error_rsc_data_out_int[19]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1350.INIT = 4'h8;
    LUT2 ix10394z1349 (.O (nx10394z28), .I0 (
         p_nbus_image_error_rsc_data_out_int[20]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1349.INIT = 4'h8;
    LUT2 ix10394z1348 (.O (nx10394z27), .I0 (
         p_nbus_image_error_rsc_data_out_int[21]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1348.INIT = 4'h8;
    LUT5 ix10394z1337 (.O (nx10394z25), .I0 (
         p_nbus_image_error_rsc_data_out_int[15]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx56642z2), .I4 (nx10394z26)) ;
         defparam ix10394z1337.INIT = 32'hECA0FFFF;
    LUT4 ix10394z3250 (.O (nx10394z26), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[8]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z10)) ;
         defparam ix10394z3250.INIT = 16'h0777;
    LUT5 ix10394z1335 (.O (nx10394z23), .I0 (
         p_nbus_image_error_rsc_data_out_int[16]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx57639z2), .I4 (nx10394z24)) ;
         defparam ix10394z1335.INIT = 32'hECA0FFFF;
    LUT4 ix10394z3248 (.O (nx10394z24), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z9)) ;
         defparam ix10394z3248.INIT = 16'h0777;
    LUT5 ix10394z1333 (.O (nx10394z21), .I0 (
         p_nbus_image_error_rsc_data_out_int[22]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx11510z4), .I4 (nx10394z22)) ;
         defparam ix10394z1333.INIT = 32'hECA0FFFF;
    LUT2 ix10394z1363 (.O (nx10394z41), .I0 (
         p_nbus_image_error_rsc_data_out_int[22]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1363.INIT = 4'h8;
    LUT4 ix10394z3246 (.O (nx10394z22), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[0]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z8)) ;
         defparam ix10394z3246.INIT = 16'h0777;
    LUT5 ix10394z1331 (.O (nx10394z19), .I0 (
         p_nbus_image_error_rsc_data_out_int[17]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx13034z3), .I4 (nx10394z20)) ;
         defparam ix10394z1331.INIT = 32'hECA0FFFF;
    LUT4 ix10394z3244 (.O (nx10394z20), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[1]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z7)) ;
         defparam ix10394z3244.INIT = 16'h0777;
    LUT5 ix10394z1329 (.O (nx10394z17), .I0 (
         p_nbus_image_error_rsc_data_out_int[18]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx12037z2), .I4 (nx10394z18)) ;
         defparam ix10394z1329.INIT = 32'hECA0FFFF;
    LUT4 ix10394z3242 (.O (nx10394z18), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[2]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z6)) ;
         defparam ix10394z3242.INIT = 16'h0777;
    LUT5 ix10394z1327 (.O (nx10394z15), .I0 (
         p_nbus_image_error_rsc_data_out_int[23]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx11040z2), .I4 (nx10394z16)) ;
         defparam ix10394z1327.INIT = 32'hECA0FFFF;
    LUT2 ix10394z1359 (.O (nx10394z38), .I0 (
         p_nbus_image_error_rsc_data_out_int[23]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1359.INIT = 4'h8;
    LUT4 ix10394z3240 (.O (nx10394z16), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z5)) ;
         defparam ix10394z3240.INIT = 16'h0777;
    LUT5 ix10394z1325 (.O (nx10394z13), .I0 (
         p_nbus_image_error_rsc_data_out_int[24]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx10043z2), .I4 (nx10394z14)) ;
         defparam ix10394z1325.INIT = 32'hECA0FFFF;
    LUT2 ix10394z1358 (.O (nx10394z37), .I0 (
         p_nbus_image_error_rsc_data_out_int[24]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1358.INIT = 4'h8;
    LUT4 ix10394z3238 (.O (nx10394z14), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z4)) ;
         defparam ix10394z3238.INIT = 16'h0777;
    LUT5 ix10394z1323 (.O (nx10394z11), .I0 (
         p_nbus_image_error_rsc_data_out_int[25]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx9046z2), .I4 (nx10394z12)) ;
         defparam ix10394z1323.INIT = 32'hECA0FFFF;
    LUT2 ix10394z1357 (.O (nx10394z36), .I0 (
         p_nbus_image_error_rsc_data_out_int[25]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1357.INIT = 4'h8;
    LUT4 ix10394z3236 (.O (nx10394z12), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z3)) ;
         defparam ix10394z3236.INIT = 16'h0777;
    LUT5 ix10394z1321 (.O (nx10394z9), .I0 (
         p_nbus_image_error_rsc_data_out_int[26]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(8)  ), .I3 (nx8049z2), .I4 (nx10394z10)) ;
         defparam ix10394z1321.INIT = 32'hECA0FFFF;
    LUT2 ix10394z1356 (.O (nx10394z35), .I0 (
         p_nbus_image_error_rsc_data_out_int[26]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1356.INIT = 4'h8;
    LUT4 ix10394z3234 (.O (nx10394z10), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[6]), .I2 (\p_for_for_mux1h_2_nl(1)  
         ), .I3 (nx4943z2)) ;
         defparam ix10394z3234.INIT = 16'h0777;
    LUT5 ix10394z5417 (.O (nx10394z8), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (p_nbus_image_error_rsc_data_out_int[27]), .I3 (
         \fsm_output(8)  ), .I4 (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[22])) ;
         defparam ix10394z5417.INIT = 32'h10111000;
    LUT2 ix10394z1355 (.O (nx10394z34), .I0 (
         p_nbus_image_error_rsc_data_out_int[27]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1355.INIT = 4'h8;
    LUT5 ix10394z5416 (.O (nx10394z7), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (p_nbus_image_error_rsc_data_out_int[28]), .I3 (
         \fsm_output(8)  ), .I4 (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[21])) ;
         defparam ix10394z5416.INIT = 32'h10111000;
    LUT2 ix10394z1354 (.O (nx10394z33), .I0 (
         p_nbus_image_error_rsc_data_out_int[28]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1354.INIT = 4'h8;
    LUT5 ix10394z5415 (.O (nx10394z6), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (p_nbus_image_error_rsc_data_out_int[29]), .I3 (
         \fsm_output(8)  ), .I4 (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[20])) ;
         defparam ix10394z5415.INIT = 32'h10111000;
    LUT2 ix10394z1353 (.O (nx10394z32), .I0 (
         p_nbus_image_error_rsc_data_out_int[29]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1353.INIT = 4'h8;
    LUT5 ix10394z5414 (.O (nx10394z5), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (p_nbus_image_error_rsc_data_out_int[30]), .I3 (
         \fsm_output(8)  ), .I4 (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[19])) ;
         defparam ix10394z5414.INIT = 32'h10111000;
    LUT2 ix10394z1352 (.O (nx10394z31), .I0 (
         p_nbus_image_error_rsc_data_out_int[30]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1352.INIT = 4'h8;
    LUT5 ix10394z5413 (.O (nx10394z4), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (p_nbus_image_error_rsc_data_out_int[31]), .I3 (
         \fsm_output(8)  ), .I4 (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[18])) ;
         defparam ix10394z5413.INIT = 32'h10111000;
    LUT2 ix10394z1351 (.O (nx10394z30), .I0 (
         p_nbus_image_error_rsc_data_out_int[31]), .I1 (\fsm_output(8)  )) ;
         defparam ix10394z1351.INIT = 4'h8;
    LUT4 ix10394z1318 (.O (nx10394z3), .I0 (
         p_nbus_image_error_rsc_data_out_int[19]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix10394z1318.INIT = 16'h0002;
    LUT4 ix10394z1317 (.O (nx10394z2), .I0 (
         p_nbus_image_error_rsc_data_out_int[20]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix10394z1317.INIT = 16'h0002;
    LUT4 ix10394z1316 (.O (nx10394z1), .I0 (
         p_nbus_image_error_rsc_data_out_int[21]), .I1 (\p_fsm_output(10)  ), .I2 (
         \fsm_output(1)  ), .I3 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix10394z1316.INIT = 16'h0002;
    LUT3 ix23312z1354 (.O (nx23312z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[15]), .I2 (\z_out(13)  
         )) ;
         defparam ix23312z1354.INIT = 8'h28;
    LUT4 ix23311z32874 (.O (nx23311z2), .I0 (
         main_core_inst_reconstruction_error_for_l_sva_3[16]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (\z_out(12)  ), .I3 (
         main_core_inst_for_for_else_acc_itm_2[1])) ;
         defparam ix23311z32874.INIT = 16'h7B48;
    LUT3 ix38388z1498 (.O (nx38388z1), .I0 (\z_out(12)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         main_core_inst_for_for_else_acc_itm_2[1])) ;
         defparam ix38388z1498.INIT = 8'hB8;
    LUT4 ix23310z32874 (.O (nx23310z2), .I0 (
         main_core_inst_reconstruction_error_for_l_sva_3[17]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (\z_out(11)  ), .I3 (
         main_core_inst_for_for_else_acc_itm_2[2])) ;
         defparam ix23310z32874.INIT = 16'h7B48;
    LUT3 ix38387z1498 (.O (nx38387z1), .I0 (\z_out(11)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         main_core_inst_for_for_else_acc_itm_2[2])) ;
         defparam ix38387z1498.INIT = 8'hB8;
    LUT4 ix23309z32874 (.O (nx23309z2), .I0 (
         main_core_inst_reconstruction_error_for_l_sva_3[18]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (\z_out(10)  ), .I3 (
         main_core_inst_for_for_else_acc_itm_2[3])) ;
         defparam ix23309z32874.INIT = 16'h7B48;
    LUT3 ix38386z1498 (.O (nx38386z1), .I0 (\z_out(10)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         main_core_inst_for_for_else_acc_itm_2[3])) ;
         defparam ix38386z1498.INIT = 8'hB8;
    LUT4 ix33887z32874 (.O (nx33887z2), .I0 (
         main_core_inst_reconstruction_error_for_l_sva_3[19]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (\z_out(9)  ), .I3 (
         main_core_inst_for_for_else_acc_itm_2[4])) ;
         defparam ix33887z32874.INIT = 16'h7B48;
    LUT3 ix26274z1498 (.O (nx26274z1), .I0 (\z_out(9)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         main_core_inst_for_for_else_acc_itm_2[4])) ;
         defparam ix26274z1498.INIT = 8'hB8;
    LUT3 ix33888z1354 (.O (nx33888z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[20]), .I2 (\p_z_out(8)  
         )) ;
         defparam ix33888z1354.INIT = 8'h28;
    LUT3 ix33889z1354 (.O (nx33889z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[21]), .I2 (\p_z_out(7)  
         )) ;
         defparam ix33889z1354.INIT = 8'h28;
    LUT3 ix33890z1354 (.O (nx33890z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[22]), .I2 (\p_z_out(6)  
         )) ;
         defparam ix33890z1354.INIT = 8'h28;
    LUT3 ix33891z1354 (.O (nx33891z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[23]), .I2 (\p_z_out(5)  
         )) ;
         defparam ix33891z1354.INIT = 8'h28;
    LUT3 ix33892z1354 (.O (nx33892z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[24]), .I2 (\p_z_out(4)  
         )) ;
         defparam ix33892z1354.INIT = 8'h28;
    LUT3 ix33893z1354 (.O (nx33893z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[25]), .I2 (\p_z_out(3)  
         )) ;
         defparam ix33893z1354.INIT = 8'h28;
    LUT3 ix33894z1354 (.O (nx33894z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[26]), .I2 (\p_z_out(2)  
         )) ;
         defparam ix33894z1354.INIT = 8'h28;
    LUT3 ix33895z1354 (.O (nx33895z2), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[27]), .I2 (\p_z_out(1)  
         )) ;
         defparam ix33895z1354.INIT = 8'h28;
    LUT3 ix33896z1354 (.O (nx33896z1), .I0 (\p_for_for_mux1h_2_nl(1)  ), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[28]), .I2 (\p_z_out(0)  
         )) ;
         defparam ix33896z1354.INIT = 8'h28;
    LUT5 ix7977z2083 (.O (nx7977z6), .I0 (nx7977z7), .I1 (nx7975z3), .I2 (
         nx7976z3), .I3 (nx7977z5), .I4 (nx7977z3)) ;
         defparam ix7977z2083.INIT = 32'hFD0202FD;
    LUT6 ix7977z1316 (.O (nx7977z2), .I0 (nx7972z2), .I1 (nx7973z3), .I2 (
         nx7975z6), .I3 (nx7975z3), .I4 (nx7976z3), .I5 (nx7977z3)) ;
         defparam ix7977z1316.INIT = 64'hFFFFFFFD00000002;
    LUT6 ix7977z18791 (.O (nx7977z3), .I0 (\fsm_output(5)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[6]), .I2 (nx7976z4), .I3 (nx7976z5)
         , .I4 (nx7977z4), .I5 (nx7977z5)) ;
         defparam ix7977z18791.INIT = 64'hEE4EEEEE44E44444;
    (* HLUTNM = "LUT62_1_27" *)
    LUT5 ix7977z53745 (.O (nx7977z5), .I0 (\for_1_i_7_0_sva_4(4)  ), .I1 (
         nx63944z3), .I2 (nx56495z7), .I3 (nx64941z4), .I4 (nx1399z3)) ;
         defparam ix7977z53745.INIT = 32'h6CCCCCCC;
    LUT6 ix7976z1315 (.O (nx7976z6), .I0 (nx7972z2), .I1 (nx7973z3), .I2 (
         nx7975z6), .I3 (nx7975z3), .I4 (nx7976z5), .I5 (nx7976z3)) ;
         defparam ix7976z1315.INIT = 64'hFFFD00020002FFFD;
    LUT5 ix7976z1316 (.O (nx7976z2), .I0 (nx7972z2), .I1 (nx7973z3), .I2 (
         nx7975z6), .I3 (nx7975z3), .I4 (nx7976z3)) ;
         defparam ix7976z1316.INIT = 32'hFFFD0002;
    LUT6 ix7976z18951 (.O (nx7976z3), .I0 (\fsm_output(5)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[5]), .I2 (nx7976z4), .I3 (nx7974z5)
         , .I4 (nx7975z8), .I5 (nx7976z5)) ;
         defparam ix7976z18951.INIT = 64'hEEEEEE4E444444E4;
    (* HLUTNM = "LUT62_1_40" *)
    LUT3 ix7977z1445 (.O (nx7977z4), .I0 (\for_1_i_7_0_sva_4(4)  ), .I1 (
         nx1399z3), .I2 (nx64941z4)) ;
         defparam ix7977z1445.INIT = 8'h81;
    (* HLUTNM = "LUT62_1_27" *)
    LUT4 ix7976z29169 (.O (nx7976z5), .I0 (\for_1_i_7_0_sva_4(4)  ), .I1 (
         nx56495z7), .I2 (nx64941z4), .I3 (nx1399z3)) ;
         defparam ix7976z29169.INIT = 16'h6CCC;
    LUT5 ix7975z2082 (.O (nx7975z5), .I0 (nx7972z2), .I1 (nx7973z3), .I2 (
         nx7975z6), .I3 (nx7975z8), .I4 (nx7975z3)) ;
         defparam ix7975z2082.INIT = 32'hFD0202FD;
    LUT6 ix7975z1330 (.O (nx7975z2), .I0 (\fsm_output(5)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (nx7972z2), .I3 (nx7973z3)
         , .I4 (nx7974z3), .I5 (nx7975z3)) ;
         defparam ix7975z1330.INIT = 64'hFF4FFFEF00B00010;
    LUT6 ix7975z62311 (.O (nx7975z3), .I0 (\fsm_output(5)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I2 (\for_1_i_7_0_sva_4(4)  ), 
         .I3 (nx64941z4), .I4 (nx1399z3), .I5 (nx7975z4)) ;
         defparam ix7975z62311.INIT = 64'hE44EEE444EE4EE44;
    (* HLUTNM = "LUT62_1_40" *)
    LUT3 ix7975z1428 (.O (nx7975z8), .I0 (\for_1_i_7_0_sva_4(4)  ), .I1 (
         nx64941z4), .I2 (nx1399z3)) ;
         defparam ix7975z1428.INIT = 8'h6C;
    LUT6 ix7974z5893 (.O (nx7974z4), .I0 (\fsm_output(5)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (nx7972z2), .I3 (nx7973z3)
         , .I4 (nx7974z5), .I5 (nx7974z3)) ;
         defparam ix7974z5893.INIT = 64'h44B4BB4BEE1E11E1;
    LUT5 ix7974z62272 (.O (nx7974z2), .I0 (\fsm_output(5)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (nx7972z2), .I3 (nx7973z3)
         , .I4 (nx7974z3)) ;
         defparam ix7974z62272.INIT = 32'h44B4EE1E;
    LUT5 ix7977z1335 (.O (nx7977z7), .I0 (\fsm_output(5)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (nx7972z2), .I3 (nx7973z3)
         , .I4 (nx7974z3)) ;
         defparam ix7977z1335.INIT = 32'h00B00010;
    LUT6 ix7975z342 (.O (nx7975z6), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         \fsm_output(5)  ), .I2 (main_core_inst_for_for_j_8_0_sva_3[3]), .I3 (
         \for_1_i_7_0_sva_4(4)  ), .I4 (nx1399z3), .I5 (nx7975z7)) ;
         defparam ix7975z342.INIT = 64'hFC30FC3074B8FC30;
    (* HLUTNM = "LUT62_1_3" *)
    LUT5 ix7974z1570 (.O (nx7974z3), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \for_1_i_7_0_sva_4(4)  ), .I4 (nx1399z3)) ;
         defparam ix7974z1570.INIT = 32'hA85700FF;
    (* HLUTNM = "LUT62_1_3" *)
    LUT5 ix7975z1403 (.O (nx7975z4), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \for_1_i_7_0_sva_4(4)  ), .I4 (nx1399z3)) ;
         defparam ix7975z1403.INIT = 32'h57000057;
    (* HLUTNM = "LUT62_1_43" *)
    LUT2 ix7974z1323 (.O (nx7974z5), .I0 (\for_1_i_7_0_sva_4(4)  ), .I1 (
         nx1399z3)) ;
         defparam ix7974z1323.INIT = 4'h6;
    LUT6 ix7973z44833 (.O (nx7973z2), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \fsm_output(5)  ), .I4 (main_core_inst_for_for_j_8_0_sva_3[1]), .I5 (
         nx7973z3)) ;
         defparam ix7973z44833.INIT = 64'h56FF5600A900A9FF;
    LUT6 ix7973z44323 (.O (nx7973z3), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \fsm_output(5)  ), .I4 (main_core_inst_for_for_j_8_0_sva_3[2]), .I5 (
         nx1399z3)) ;
         defparam ix7973z44323.INIT = 64'h57FF5700A8FFA800;
    (* HLUTNM = "LUT62_1_56" *)
    LUT4 ix7976z23588 (.O (nx7976z4), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         nx1399z3)) ;
         defparam ix7976z23588.INIT = 16'h5700;
    LUT5 ix7972z461 (.O (nx7972z3), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \fsm_output(5)  ), .I4 (main_core_inst_for_for_j_8_0_sva_3[1])) ;
         defparam ix7972z461.INIT = 32'hFC55FCAA;
    LUT5 ix7972z44833 (.O (nx7972z2), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         p_nbus_depth_rsc_addr_1_0[1]), .I2 (p_nbus_depth_rsc_addr_1_0[0]), .I3 (
         \fsm_output(5)  ), .I4 (main_core_inst_for_for_j_8_0_sva_3[1])) ;
         defparam ix7972z44833.INIT = 32'hA900A9FF;
    LUT2 ix7971z1324 (.O (nx7971z1), .I0 (p_nbus_depth_rsc_addr_1_0[1]), .I1 (
         p_nbus_depth_rsc_addr_1_0[0])) ;
         defparam ix7971z1324.INIT = 4'h9;
    (* HLUTNM = "LUT62_1_41" *)
    LUT2 ix7975z1320 (.O (nx7975z7), .I0 (p_nbus_depth_rsc_addr_1_0[1]), .I1 (
         p_nbus_depth_rsc_addr_1_0[0])) ;
         defparam ix7975z1320.INIT = 4'h1;
    LUT3 ix34912z1540 (.O (nx34912z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[1]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[30])) ;
         defparam ix34912z1540.INIT = 8'hE2;
    LUT3 ix33924z1540 (.O (nx33924z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[2]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[29])) ;
         defparam ix33924z1540.INIT = 8'hE2;
    LUT3 ix33923z1540 (.O (nx33923z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[3]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[28])) ;
         defparam ix33923z1540.INIT = 8'hE2;
    LUT3 ix33922z1540 (.O (nx33922z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[4]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[27])) ;
         defparam ix33922z1540.INIT = 8'hE2;
    LUT3 ix33921z1540 (.O (nx33921z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[5]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[26])) ;
         defparam ix33921z1540.INIT = 8'hE2;
    LUT3 ix33920z1540 (.O (nx33920z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[6]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[25])) ;
         defparam ix33920z1540.INIT = 8'hE2;
    LUT3 ix33919z1540 (.O (nx33919z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[7]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[24])) ;
         defparam ix33919z1540.INIT = 8'hE2;
    LUT3 ix33918z1540 (.O (nx33918z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[8]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[23])) ;
         defparam ix33918z1540.INIT = 8'hE2;
    LUT3 ix33917z1540 (.O (nx33917z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[9]), .I1 (nx31299z1
         ), .I2 (p_nbus_image_floue_rsc_data_out_int[22])) ;
         defparam ix33917z1540.INIT = 8'hE2;
    LUT3 ix33916z1540 (.O (nx33916z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[10]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[21])) ;
         defparam ix33916z1540.INIT = 8'hE2;
    LUT3 ix33915z1540 (.O (nx33915z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[11]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[20])) ;
         defparam ix33915z1540.INIT = 8'hE2;
    LUT3 ix32927z1540 (.O (nx32927z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[12]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[19])) ;
         defparam ix32927z1540.INIT = 8'hE2;
    LUT3 ix32926z1540 (.O (nx32926z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[13]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[18])) ;
         defparam ix32926z1540.INIT = 8'hE2;
    LUT3 ix32925z1540 (.O (nx32925z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[14]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[17])) ;
         defparam ix32925z1540.INIT = 8'hE2;
    LUT3 ix32924z1540 (.O (nx32924z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[15]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[16])) ;
         defparam ix32924z1540.INIT = 8'hE2;
    LUT3 ix32923z1540 (.O (nx32923z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[16]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[15])) ;
         defparam ix32923z1540.INIT = 8'hE2;
    LUT3 ix32922z1540 (.O (nx32922z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[17]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[14])) ;
         defparam ix32922z1540.INIT = 8'hE2;
    LUT3 ix32921z1540 (.O (nx32921z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[18]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[13])) ;
         defparam ix32921z1540.INIT = 8'hE2;
    LUT3 ix32920z1540 (.O (nx32920z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[19]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[12])) ;
         defparam ix32920z1540.INIT = 8'hE2;
    LUT3 ix32919z1540 (.O (nx32919z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[20]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[11])) ;
         defparam ix32919z1540.INIT = 8'hE2;
    LUT3 ix32918z1540 (.O (nx32918z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[21]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[10])) ;
         defparam ix32918z1540.INIT = 8'hE2;
    LUT3 ix17526z1540 (.O (nx17526z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[22]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[9])) ;
         defparam ix17526z1540.INIT = 8'hE2;
    LUT3 ix17525z1540 (.O (nx17525z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[23]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[8])) ;
         defparam ix17525z1540.INIT = 8'hE2;
    LUT3 ix17524z1540 (.O (nx17524z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[24]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[7])) ;
         defparam ix17524z1540.INIT = 8'hE2;
    LUT3 ix17523z1540 (.O (nx17523z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[25]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[6])) ;
         defparam ix17523z1540.INIT = 8'hE2;
    LUT3 ix17522z1540 (.O (nx17522z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[26]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[5])) ;
         defparam ix17522z1540.INIT = 8'hE2;
    LUT3 ix17521z1540 (.O (nx17521z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[27]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[4])) ;
         defparam ix17521z1540.INIT = 8'hE2;
    LUT3 ix17520z1540 (.O (nx17520z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[28]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[3])) ;
         defparam ix17520z1540.INIT = 8'hE2;
    LUT3 ix17519z1540 (.O (nx17519z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[29]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[2])) ;
         defparam ix17519z1540.INIT = 8'hE2;
    LUT3 ix17518z1540 (.O (nx17518z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[30]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[1])) ;
         defparam ix17518z1540.INIT = 8'hE2;
    LUT3 ix17517z1540 (.O (nx17517z1), .I0 (
         main_core_inst_reconstruction_error_rec_error_lpi_6[31]), .I1 (
         nx31299z1), .I2 (p_nbus_image_floue_rsc_data_out_int[0])) ;
         defparam ix17517z1540.INIT = 8'hE2;
    LUT4 ix50036z40542 (.O (nx50036z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[5]), .I1 (nx39519z1), .I2 (
         nx39519z3), .I3 (nx21269z2)) ;
         defparam ix50036z40542.INIT = 16'h993C;
    LUT3 ix39524z1420 (.O (nx39524z3), .I0 (nx39524z2), .I1 (nx39519z3), .I2 (
         nx21269z2)) ;
         defparam ix39524z1420.INIT = 8'h69;
    LUT6 ix21269z1316 (.O (nx21269z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2]), .I1 (nx21269z3), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[4]), .I3 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[3]), .I4 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I5 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0])) ;
         defparam ix21269z1316.INIT = 64'h0000000000000001;
    LUT6 ix39524z1314 (.O (nx39524z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[4]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[3]), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2]), .I3 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I4 (nx39519z3), .I5 (
         nx23263z2)) ;
         defparam ix39524z1314.INIT = 64'hFFFD0001FFFF0000;
    LUT5 ix39523z1058 (.O (nx39523z3), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I3 (nx39519z3), .I4 (
         nx21269z3)) ;
         defparam ix39523z1058.INIT = 32'hFFFFFEFF;
    LUT5 ix22266z1316 (.O (nx22266z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I1 (nx21269z3), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I3 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[3]), .I4 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2])) ;
         defparam ix22266z1316.INIT = 32'h00000001;
    LUT6 ix39523z1315 (.O (nx39523z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[3]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2]), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I3 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I4 (nx39519z3), .I5 (
         nx21269z3)) ;
         defparam ix39523z1315.INIT = 64'hFFFF0000FFFD0001;
    LUT6 ix39522z62738 (.O (nx39522z3), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I2 (nx39519z3), .I3 (
         nx11510z4), .I4 (nx57639z2), .I5 (nx56642z2)) ;
         defparam ix39522z62738.INIT = 64'hFFEFFFEFFFEFEFEF;
    LUT5 ix39522z547 (.O (nx39522z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[2]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I2 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I3 (nx39519z3), .I4 (
         nx21269z3)) ;
         defparam ix39522z547.INIT = 32'hFF00FD01;
    LUT5 ix39521z222 (.O (nx39521z3), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I1 (nx39519z3), .I2 (
         nx11510z4), .I3 (nx57639z2), .I4 (nx56642z2)) ;
         defparam ix39521z222.INIT = 32'hFBFBFBBB;
    LUT6 ix39521z55027 (.O (nx39521z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[1]), .I1 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I2 (nx39519z3), .I3 (
         nx11510z4), .I4 (nx57639z2), .I5 (nx56642z2)) ;
         defparam ix39521z55027.INIT = 64'hF0D1F0D1F0D1D1D1;
    LUT4 ix39520z58104 (.O (nx39520z3), .I0 (nx39519z3), .I1 (nx11510z4), .I2 (
         nx57639z2), .I3 (nx56642z2)) ;
         defparam ix39520z58104.INIT = 16'hDDD5;
    LUT4 ix23263z5688 (.O (nx23263z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I1 (nx11510z4), .I2 (
         nx57639z2), .I3 (nx56642z2)) ;
         defparam ix23263z5688.INIT = 16'h1115;
    LUT5 ix39520z51831 (.O (nx39520z2), .I0 (
         main_core_inst_for_1_for_acc_7_psp_1_sva_1[0]), .I1 (nx39519z3), .I2 (
         nx11510z4), .I3 (nx57639z2), .I4 (nx56642z2)) ;
         defparam ix39520z51831.INIT = 32'hC5C5C555;
    (* HLUTNM = "LUT62_1_38" *)
    LUT3 ix21269z1484 (.O (nx21269z3), .I0 (nx11510z4), .I1 (nx57639z2), .I2 (
         nx56642z2)) ;
         defparam ix21269z1484.INIT = 8'hA8;
    LUT4 ix39519z14429 (.O (nx39519z2), .I0 (nx39519z3), .I1 (nx11510z4), .I2 (
         nx57639z2), .I3 (nx56642z2)) ;
         defparam ix39519z14429.INIT = 16'h333A;
    LUT3 ix34672z1530 (.O (nx34672z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[1]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[1])) ;
         defparam ix34672z1530.INIT = 8'hD8;
    LUT3 ix35660z1530 (.O (nx35660z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[2]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[2])) ;
         defparam ix35660z1530.INIT = 8'hD8;
    LUT3 ix35661z1530 (.O (nx35661z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[3]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[3])) ;
         defparam ix35661z1530.INIT = 8'hD8;
    LUT3 ix35662z1530 (.O (nx35662z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[4]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[4])) ;
         defparam ix35662z1530.INIT = 8'hD8;
    LUT3 ix35663z1530 (.O (nx35663z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[5]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[5])) ;
         defparam ix35663z1530.INIT = 8'hD8;
    LUT3 ix35664z1530 (.O (nx35664z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[6]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[6])) ;
         defparam ix35664z1530.INIT = 8'hD8;
    LUT3 ix35665z1530 (.O (nx35665z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[7]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[7])) ;
         defparam ix35665z1530.INIT = 8'hD8;
    LUT3 ix35666z1530 (.O (nx35666z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[8]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[8])) ;
         defparam ix35666z1530.INIT = 8'hD8;
    LUT3 ix35667z1530 (.O (nx35667z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[9]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[9])) ;
         defparam ix35667z1530.INIT = 8'hD8;
    LUT3 ix35668z1530 (.O (nx35668z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[10]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[10])) ;
         defparam ix35668z1530.INIT = 8'hD8;
    LUT3 ix35669z1530 (.O (nx35669z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[11]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[11])) ;
         defparam ix35669z1530.INIT = 8'hD8;
    LUT3 ix36657z1530 (.O (nx36657z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[12]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[12])) ;
         defparam ix36657z1530.INIT = 8'hD8;
    LUT3 ix36658z1530 (.O (nx36658z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[13]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[13])) ;
         defparam ix36658z1530.INIT = 8'hD8;
    LUT3 ix36659z1530 (.O (nx36659z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[14]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[14])) ;
         defparam ix36659z1530.INIT = 8'hD8;
    LUT3 ix36660z1530 (.O (nx36660z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[15]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[15])) ;
         defparam ix36660z1530.INIT = 8'hD8;
    LUT3 ix36661z1530 (.O (nx36661z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[16]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[16])) ;
         defparam ix36661z1530.INIT = 8'hD8;
    LUT3 ix36662z1530 (.O (nx36662z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[17]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[17])) ;
         defparam ix36662z1530.INIT = 8'hD8;
    LUT3 ix36663z1530 (.O (nx36663z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[18]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[18])) ;
         defparam ix36663z1530.INIT = 8'hD8;
    LUT3 ix36664z1530 (.O (nx36664z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[19]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[19])) ;
         defparam ix36664z1530.INIT = 8'hD8;
    LUT3 ix36665z1530 (.O (nx36665z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[20]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[20])) ;
         defparam ix36665z1530.INIT = 8'hD8;
    LUT3 ix36666z1530 (.O (nx36666z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[21]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[21])) ;
         defparam ix36666z1530.INIT = 8'hD8;
    LUT3 ix12058z1530 (.O (nx12058z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[22]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[22])) ;
         defparam ix12058z1530.INIT = 8'hD8;
    LUT3 ix12059z1530 (.O (nx12059z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[23]), .I2 (
         main_core_inst_z_out_8[0])) ;
         defparam ix12059z1530.INIT = 8'hD8;
    LUT4 ix12060z55045 (.O (nx12060z3), .I0 (nx12060z4), .I1 (\p_fsm_output(10)  
         ), .I2 (main_core_inst_reconstruction_error_rec_error_sva[24]), .I3 (
         main_core_inst_z_out_8[1])) ;
         defparam ix12060z55045.INIT = 16'hD1E2;
    LUT5 ix12060z62841 (.O (nx12060z4), .I0 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[0]), .I1 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[1]), .I2 (
         main_core_inst_z_out_2[5]), .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (
         nx12061z4)) ;
         defparam ix12060z62841.INIT = 32'hF099F055;
    LUT3 ix12060z1530 (.O (nx12060z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[24]), .I2 (
         main_core_inst_z_out_8[1])) ;
         defparam ix12060z1530.INIT = 8'hD8;
    LUT6 ix12061z21812 (.O (nx12061z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[1]), .I2 (
         main_core_inst_z_out_2[4]), .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (
         nx12061z2), .I5 (nx12061z4)) ;
         defparam ix12061z21812.INIT = 64'hAFBB5044AFEE5011;
    (* HLUTNM = "LUT62_1_44" *)
    LUT4 ix12061z34084 (.O (nx12061z4), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[4]), .I2 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[2]), .I3 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[3])) ;
         defparam ix12061z34084.INIT = 16'h8000;
    LUT3 ix12061z1530 (.O (nx12061z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[25]), .I2 (
         main_core_inst_z_out_8[2])) ;
         defparam ix12061z1530.INIT = 8'hD8;
    LUT4 ix12062z55045 (.O (nx12062z3), .I0 (nx12062z4), .I1 (\p_fsm_output(10)  
         ), .I2 (main_core_inst_reconstruction_error_rec_error_sva[26]), .I3 (
         main_core_inst_z_out_8[3])) ;
         defparam ix12062z55045.INIT = 16'hD1E2;
    LUT6 ix12062z38999 (.O (nx12062z4), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[2]), .I2 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[3]), .I3 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[4]), .I4 (
         main_core_inst_z_out_2[3]), .I5 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix12062z38999.INIT = 64'hFFFF000093339333;
    LUT3 ix12062z1530 (.O (nx12062z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[26]), .I2 (
         main_core_inst_z_out_8[3])) ;
         defparam ix12062z1530.INIT = 8'hD8;
    LUT6 ix12063z21812 (.O (nx12063z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[3]), .I2 (
         main_core_inst_z_out_2[2]), .I3 (\p_for_for_mux1h_2_nl(1)  ), .I4 (
         nx12063z2), .I5 (nx12063z4)) ;
         defparam ix12063z21812.INIT = 64'hAFBB5044AFEE5011;
    (* HLUTNM = "LUT62_1_44" *)
    LUT2 ix12063z1324 (.O (nx12063z4), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[4])) ;
         defparam ix12063z1324.INIT = 4'h8;
    LUT3 ix12063z1530 (.O (nx12063z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[27]), .I2 (
         main_core_inst_z_out_8[4])) ;
         defparam ix12063z1530.INIT = 8'hD8;
    LUT6 ix12064z9796 (.O (nx12064z3), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         \p_fsm_output(10)  ), .I2 (
         main_core_inst_for_1_for_acc_6_psp_1_sva_1[4]), .I3 (
         main_core_inst_z_out_2[1]), .I4 (\p_for_for_mux1h_2_nl(1)  ), .I5 (
         nx12064z2)) ;
         defparam ix12064z9796.INIT = 64'hCCFFDEDE33002121;
    LUT3 ix12064z1530 (.O (nx12064z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[28]), .I2 (
         main_core_inst_z_out_8[5])) ;
         defparam ix12064z1530.INIT = 8'hD8;
    LUT6 ix12065z59397 (.O (nx12065z3), .I0 (p_nbus_depth_rsc_addr_1_0[2]), .I1 (
         \p_fsm_output(10)  ), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[29]), .I3 (
         main_core_inst_z_out_2[0]), .I4 (main_core_inst_z_out_8[6]), .I5 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix12065z59397.INIT = 64'hC0F3F3C0D1D1E2E2;
    LUT3 ix12065z1530 (.O (nx12065z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[29]), .I2 (
         main_core_inst_z_out_8[6])) ;
         defparam ix12065z1530.INIT = 8'hD8;
    LUT3 ix12066z1530 (.O (nx12066z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[30]), .I2 (
         main_core_inst_z_out_8[7])) ;
         defparam ix12066z1530.INIT = 8'hD8;
    LUT3 ix12067z1530 (.O (nx12067z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[31]), .I2 (
         main_core_inst_z_out_8[8])) ;
         defparam ix12067z1530.INIT = 8'hD8;
    (* HLUTNM = "LUT62_1_55" *)
    LUT2 ix11516z1329 (.O (nx11516z3), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  )) ;
         defparam ix11516z1329.INIT = 4'hE;
    LUT3 ix11510z1568 (.O (nx11510z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \fsm_output(1)  ), .I2 (\p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix11510z1568.INIT = 8'hFE;
    LUT2 ix11512z1328 (.O (nx11512z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix11512z1328.INIT = 4'hE;
    LUT3 ix40591z1530 (.O (nx40591z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \z_out(12)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[12])) ;
         defparam ix40591z1530.INIT = 8'hD8;
    LUT3 ix55667z1530 (.O (nx55667z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \z_out(11)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[11])) ;
         defparam ix55667z1530.INIT = 8'hD8;
    LUT3 ix55666z1530 (.O (nx55666z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \z_out(10)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[10])) ;
         defparam ix55666z1530.INIT = 8'hD8;
    LUT3 ix25634z1530 (.O (nx25634z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \z_out(9)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[9])) ;
         defparam ix25634z1530.INIT = 8'hD8;
    LUT3 ix25633z1530 (.O (nx25633z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \p_z_out(8)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[8])) ;
         defparam ix25633z1530.INIT = 8'hD8;
    LUT3 ix25632z1530 (.O (nx25632z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \p_z_out(7)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[7])) ;
         defparam ix25632z1530.INIT = 8'hD8;
    LUT3 ix25631z1530 (.O (nx25631z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \p_z_out(6)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[6])) ;
         defparam ix25631z1530.INIT = 8'hD8;
    LUT3 ix25630z1530 (.O (nx25630z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \p_z_out(5)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[5])) ;
         defparam ix25630z1530.INIT = 8'hD8;
    LUT3 ix25629z1530 (.O (nx25629z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \p_z_out(4)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[4])) ;
         defparam ix25629z1530.INIT = 8'hD8;
    LUT3 ix25628z1530 (.O (nx25628z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \p_z_out(3)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[3])) ;
         defparam ix25628z1530.INIT = 8'hD8;
    LUT3 ix25627z1530 (.O (nx25627z2), .I0 (\p_fsm_output(10)  ), .I1 (
         \p_z_out(2)  ), .I2 (main_core_inst_for_for_else_mul_2_nl[2])) ;
         defparam ix25627z1530.INIT = 8'hD8;
    LUT3 ix25626z1542 (.O (nx25626z2), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I2 (\p_z_out(1)  )) ;
         defparam ix25626z1542.INIT = 8'hE4;
    LUT3 ix25625z1542 (.O (nx25625z1), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_for_for_j_8_0_sva_3[8]), .I2 (\p_z_out(0)  )) ;
         defparam ix25625z1542.INIT = 8'hE4;
    LUT3 ix4943z1498 (.O (nx4943z1), .I0 (
         main_core_inst_reconstruction_error_for_for_c_sva_31_9_2[0]), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         main_core_inst_reconstruction_error_for_l_sva_3[0])) ;
         defparam ix4943z1498.INIT = 8'hB8;
    (* HLUTNM = "LUT62_1_100" *)
    LUT2 ix57058z1327 (.O (px1827), .I0 (\fsm_output(1)  ), .I1 (nx6053z1)) ;
         defparam ix57058z1327.INIT = 4'hD;
    LUT2 ix57057z1322 (.O (px1828), .I0 (main_core_inst_z_out_6[31]), .I1 (
         nx31299z1)) ;
         defparam ix57057z1322.INIT = 4'h8;
    LUT2 ix57056z1322 (.O (px1829), .I0 (main_core_inst_z_out_6[30]), .I1 (
         nx31299z1)) ;
         defparam ix57056z1322.INIT = 4'h8;
    LUT2 ix56068z1322 (.O (px1830), .I0 (main_core_inst_z_out_6[29]), .I1 (
         nx31299z1)) ;
         defparam ix56068z1322.INIT = 4'h8;
    LUT2 ix56067z1322 (.O (px1831), .I0 (main_core_inst_z_out_6[28]), .I1 (
         nx31299z1)) ;
         defparam ix56067z1322.INIT = 4'h8;
    LUT2 ix56066z1322 (.O (px1832), .I0 (main_core_inst_z_out_6[27]), .I1 (
         nx31299z1)) ;
         defparam ix56066z1322.INIT = 4'h8;
    LUT2 ix56065z1322 (.O (px1833), .I0 (main_core_inst_z_out_6[26]), .I1 (
         nx31299z1)) ;
         defparam ix56065z1322.INIT = 4'h8;
    LUT2 ix56064z1322 (.O (px1834), .I0 (main_core_inst_z_out_6[25]), .I1 (
         nx31299z1)) ;
         defparam ix56064z1322.INIT = 4'h8;
    LUT2 ix56063z1322 (.O (px1835), .I0 (main_core_inst_z_out_6[24]), .I1 (
         nx31299z1)) ;
         defparam ix56063z1322.INIT = 4'h8;
    LUT2 ix56062z1322 (.O (px1836), .I0 (main_core_inst_z_out_6[23]), .I1 (
         nx31299z1)) ;
         defparam ix56062z1322.INIT = 4'h8;
    LUT2 ix56061z1322 (.O (px1837), .I0 (main_core_inst_z_out_6[22]), .I1 (
         nx31299z1)) ;
         defparam ix56061z1322.INIT = 4'h8;
    LUT2 ix56060z1322 (.O (px1838), .I0 (main_core_inst_z_out_6[21]), .I1 (
         nx31299z1)) ;
         defparam ix56060z1322.INIT = 4'h8;
    LUT2 ix56059z1322 (.O (px1839), .I0 (main_core_inst_z_out_6[20]), .I1 (
         nx31299z1)) ;
         defparam ix56059z1322.INIT = 4'h8;
    LUT2 ix55071z1322 (.O (px1840), .I0 (main_core_inst_z_out_6[19]), .I1 (
         nx31299z1)) ;
         defparam ix55071z1322.INIT = 4'h8;
    LUT2 ix55070z1322 (.O (px1841), .I0 (main_core_inst_z_out_6[18]), .I1 (
         nx31299z1)) ;
         defparam ix55070z1322.INIT = 4'h8;
    LUT2 ix55069z1322 (.O (px1842), .I0 (main_core_inst_z_out_6[17]), .I1 (
         nx31299z1)) ;
         defparam ix55069z1322.INIT = 4'h8;
    LUT2 ix55068z1322 (.O (px1843), .I0 (main_core_inst_z_out_6[16]), .I1 (
         nx31299z1)) ;
         defparam ix55068z1322.INIT = 4'h8;
    LUT2 ix55067z1322 (.O (px1844), .I0 (main_core_inst_z_out_6[15]), .I1 (
         nx31299z1)) ;
         defparam ix55067z1322.INIT = 4'h8;
    LUT2 ix55066z1322 (.O (px1845), .I0 (main_core_inst_z_out_6[14]), .I1 (
         nx31299z1)) ;
         defparam ix55066z1322.INIT = 4'h8;
    LUT2 ix55065z1322 (.O (px1846), .I0 (main_core_inst_z_out_6[13]), .I1 (
         nx31299z1)) ;
         defparam ix55065z1322.INIT = 4'h8;
    LUT2 ix55064z1322 (.O (px1847), .I0 (main_core_inst_z_out_6[12]), .I1 (
         nx31299z1)) ;
         defparam ix55064z1322.INIT = 4'h8;
    LUT2 ix55063z1322 (.O (px1848), .I0 (main_core_inst_z_out_6[11]), .I1 (
         nx31299z1)) ;
         defparam ix55063z1322.INIT = 4'h8;
    LUT2 ix55062z1322 (.O (px1849), .I0 (main_core_inst_z_out_6[10]), .I1 (
         nx31299z1)) ;
         defparam ix55062z1322.INIT = 4'h8;
    LUT2 ix54074z1322 (.O (px1850), .I0 (main_core_inst_z_out_6[9]), .I1 (
         nx31299z1)) ;
         defparam ix54074z1322.INIT = 4'h8;
    LUT2 ix54073z1322 (.O (px1851), .I0 (main_core_inst_z_out_6[8]), .I1 (
         nx31299z1)) ;
         defparam ix54073z1322.INIT = 4'h8;
    LUT2 ix54072z1322 (.O (px1852), .I0 (main_core_inst_z_out_6[7]), .I1 (
         nx31299z1)) ;
         defparam ix54072z1322.INIT = 4'h8;
    LUT2 ix54071z1322 (.O (px1853), .I0 (main_core_inst_z_out_6[6]), .I1 (
         nx31299z1)) ;
         defparam ix54071z1322.INIT = 4'h8;
    LUT2 ix54070z1322 (.O (px1854), .I0 (main_core_inst_z_out_6[5]), .I1 (
         nx31299z1)) ;
         defparam ix54070z1322.INIT = 4'h8;
    LUT2 ix54069z1322 (.O (px1855), .I0 (main_core_inst_z_out_6[4]), .I1 (
         nx31299z1)) ;
         defparam ix54069z1322.INIT = 4'h8;
    LUT2 ix54068z1322 (.O (px1856), .I0 (main_core_inst_z_out_6[3]), .I1 (
         nx31299z1)) ;
         defparam ix54068z1322.INIT = 4'h8;
    LUT2 ix54067z1322 (.O (px1857), .I0 (main_core_inst_z_out_6[2]), .I1 (
         nx31299z1)) ;
         defparam ix54067z1322.INIT = 4'h8;
    LUT2 ix54066z1322 (.O (px1858), .I0 (main_core_inst_z_out_6[1]), .I1 (
         nx31299z1)) ;
         defparam ix54066z1322.INIT = 4'h8;
    LUT2 ix54065z1322 (.O (px1859), .I0 (main_core_inst_z_out_6[0]), .I1 (
         nx31299z1)) ;
         defparam ix54065z1322.INIT = 4'h8;
    LUT5 ix53077z1218 (.O (px1860), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[0]), .I2 (\z_out(13)  ), .I3 (
         image_error_mux1h_nl_0n0s3), .I4 (nx31299z1)) ;
         defparam ix53077z1218.INIT = 32'hFFECFFA0;
    LUT2 ix53076z1318 (.O (px1861), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_image_error_mux_nl[3])) ;
         defparam ix53076z1318.INIT = 4'h4;
    LUT2 ix53075z1318 (.O (px1862), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_image_error_mux_nl[2])) ;
         defparam ix53075z1318.INIT = 4'h4;
    LUT2 ix53074z1318 (.O (px1863), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_image_error_mux_nl[1])) ;
         defparam ix53074z1318.INIT = 4'h4;
    LUT2 ix53073z1318 (.O (px1864), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_image_error_mux_nl[0])) ;
         defparam ix53073z1318.INIT = 4'h4;
    LUT5 ix53072z1218 (.O (px1865), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[5]), .I2 (
         main_core_inst_for_for_if_acc_nl[8]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[8]), .I4 (nx31299z1)) ;
         defparam ix53072z1218.INIT = 32'hFFECFFA0;
    LUT5 ix53071z1218 (.O (px1866), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[6]), .I2 (
         main_core_inst_for_for_if_acc_nl[7]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[7]), .I4 (nx31299z1)) ;
         defparam ix53071z1218.INIT = 32'hFFECFFA0;
    LUT5 ix53070z1218 (.O (px1867), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[7]), .I2 (
         main_core_inst_for_for_if_acc_nl[6]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[6]), .I4 (nx31299z1)) ;
         defparam ix53070z1218.INIT = 32'hFFECFFA0;
    LUT5 ix53069z1218 (.O (px1868), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[8]), .I2 (
         main_core_inst_for_for_if_acc_nl[5]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[5]), .I4 (nx31299z1)) ;
         defparam ix53069z1218.INIT = 32'hFFECFFA0;
    LUT5 ix53068z1218 (.O (px1869), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[9]), .I2 (
         main_core_inst_for_for_if_acc_nl[4]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[4]), .I4 (nx31299z1)) ;
         defparam ix53068z1218.INIT = 32'hFFECFFA0;
    LUT5 ix52080z1218 (.O (px1870), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[10]), .I2 (
         main_core_inst_for_for_if_acc_nl[3]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[3]), .I4 (nx31299z1)) ;
         defparam ix52080z1218.INIT = 32'hFFECFFA0;
    LUT5 ix52079z1218 (.O (px1871), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[11]), .I2 (
         main_core_inst_for_for_if_acc_nl[2]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[2]), .I4 (nx31299z1)) ;
         defparam ix52079z1218.INIT = 32'hFFECFFA0;
    LUT5 ix52078z1218 (.O (px1872), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[12]), .I2 (
         main_core_inst_for_for_if_acc_nl[1]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[1]), .I4 (nx31299z1)) ;
         defparam ix52078z1218.INIT = 32'hFFECFFA0;
    LUT5 ix52077z1218 (.O (px1873), .I0 (\fsm_output(1)  ), .I1 (
         main_core_inst_for_for_else_acc_itm_2[13]), .I2 (
         main_core_inst_for_for_if_acc_nl[0]), .I3 (
         main_core_inst_image_error_mux1h_2_nl_0n0s3[0]), .I4 (nx31299z1)) ;
         defparam ix52077z1218.INIT = 32'hFFECFFA0;
    LUT3 ix52076z1516 (.O (px1874), .I0 (p_nbus_image_net_rsc_addr_1_0[13]), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[29]), .I2 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix52076z1516.INIT = 8'hCA;
    (* HLUTNM = "LUT62_1_77" *)
    LUT3 ix52075z1516 (.O (px1875), .I0 (p_nbus_image_net_rsc_addr_1_0[14]), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[30]), .I2 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix52075z1516.INIT = 8'hCA;
    (* HLUTNM = "LUT62_1_77" *)
    LUT3 ix52074z1516 (.O (px1876), .I0 (p_nbus_image_net_rsc_addr_1_0[15]), .I1 (
         main_core_inst_reconstruction_error_for_l_sva_3[31]), .I2 (
         \p_for_for_mux1h_2_nl(1)  )) ;
         defparam ix52074z1516.INIT = 8'hCA;
    (* HLUTNM = "LUT62_1_55" *)
    LUT4 ix52073z19185 (.O (px1877), .I0 (\fsm_output(1)  ), .I1 (
         for_for_if_for_for_if_and_itm_1), .I2 (nx31299z1), .I3 (nx6053z1)) ;
         defparam ix52073z19185.INIT = 16'h45CF;
    LUT6 ix6053z23158 (.O (nx6053z1), .I0 (nx52183z2), .I1 (nx6053z2), .I2 (
         nx6053z3), .I3 (nx6053z4), .I4 (nx6053z5), .I5 (nx6053z6)) ;
         defparam ix6053z23158.INIT = 64'hFFFCFFFCFFFC5554;
    LUT6 ix6053z44496 (.O (nx6053z6), .I0 (main_core_inst_for_for_j_8_0_sva_3[6]
         ), .I1 (main_core_inst_for_for_j_8_0_sva_3[5]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[4]), .I3 (
         main_core_inst_for_for_j_8_0_sva_3[3]), .I4 (
         main_core_inst_for_for_j_8_0_sva_3[2]), .I5 (
         main_core_inst_for_for_j_8_0_sva_3[1])) ;
         defparam ix6053z44496.INIT = 64'hAAA8A8A8A8A8A8A8;
    LUT6 ix6053z1319 (.O (nx6053z5), .I0 (main_core_inst_for_for_j_8_0_sva_3[6])
         , .I1 (main_core_inst_for_for_j_8_0_sva_3[3]), .I2 (
         main_core_inst_for_for_j_8_0_sva_3[2]), .I3 (
         main_core_inst_for_for_j_8_0_sva_3[0]), .I4 (
         main_core_inst_for_for_j_8_0_sva_3[7]), .I5 (
         main_core_inst_for_for_j_8_0_sva_3[8])) ;
         defparam ix6053z1319.INIT = 64'h8000800080000000;
    LUT5 ix6053z1323 (.O (nx6053z4), .I0 (p_nbus_image_net_rsc_addr_1_0[13]), .I1 (
         p_nbus_image_net_rsc_addr_1_0[14]), .I2 (\for_i_7_0_sva_3(7)  ), .I3 (
         \for_i_7_0_sva_3(6)  ), .I4 (\for_i_7_0_sva_3(4)  )) ;
         defparam ix6053z1323.INIT = 32'hE0000000;
    LUT5 ix6053z1317 (.O (nx6053z3), .I0 (\for_i_7_0_sva_3(7)  ), .I1 (
         \for_i_7_0_sva_3(6)  ), .I2 (\for_i_7_0_sva_3(5)  ), .I3 (
         \for_i_7_0_sva_3(4)  ), .I4 (\for_i_7_0_sva_3(3)  )) ;
         defparam ix6053z1317.INIT = 32'h00000001;
    LUT6 ix6053z50467 (.O (nx6053z2), .I0 (p_nbus_image_net_rsc_addr_1_0[15]), .I1 (
         \for_i_7_0_sva_3(7)  ), .I2 (\for_i_7_0_sva_3(6)  ), .I3 (
         \for_i_7_0_sva_3(5)  ), .I4 (\for_i_7_0_sva_3(4)  ), .I5 (
         \for_i_7_0_sva_3(3)  )) ;
         defparam ix6053z50467.INIT = 64'hC0C0C000C080C000;
    (* HLUTNM = "LUT62_1_4" *)
    LUT4 ix51079z52718 (.O (px1884), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I3 (
         nx34290z2)) ;
         defparam ix51079z52718.INIT = 16'hC8CC;
    LUT5 ix51078z62994 (.O (px1885), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[1]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix51078z62994.INIT = 32'hD080F0F0;
    LUT5 ix51077z62994 (.O (px1886), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[2]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix51077z62994.INIT = 32'hD080F0F0;
    LUT5 ix51076z62994 (.O (px1887), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[3]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix51076z62994.INIT = 32'hD080F0F0;
    LUT5 ix51075z62994 (.O (px1888), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[4]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix51075z62994.INIT = 32'hD080F0F0;
    LUT5 ix51074z62994 (.O (px1889), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[5]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix51074z62994.INIT = 32'hD080F0F0;
    LUT5 ix50086z62994 (.O (px1890), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[6]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50086z62994.INIT = 32'hD080F0F0;
    LUT5 ix50085z62994 (.O (px1891), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[7]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50085z62994.INIT = 32'hD080F0F0;
    LUT5 ix50084z62994 (.O (px1892), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[8]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50084z62994.INIT = 32'hD080F0F0;
    LUT5 ix50083z62994 (.O (px1893), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[9]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50083z62994.INIT = 32'hD080F0F0;
    LUT5 ix50082z62994 (.O (px1894), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[10]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50082z62994.INIT = 32'hD080F0F0;
    LUT5 ix50081z62994 (.O (px1895), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[11]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50081z62994.INIT = 32'hD080F0F0;
    LUT5 ix50080z62994 (.O (px1896), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[12]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50080z62994.INIT = 32'hD080F0F0;
    LUT5 ix50079z62994 (.O (px1897), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[13]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50079z62994.INIT = 32'hD080F0F0;
    LUT5 ix50078z62994 (.O (px1898), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[14]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50078z62994.INIT = 32'hD080F0F0;
    LUT5 ix50077z62994 (.O (px1899), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[15]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix50077z62994.INIT = 32'hD080F0F0;
    LUT5 ix48090z62994 (.O (px1900), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[16]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48090z62994.INIT = 32'hD080F0F0;
    LUT5 ix48089z62994 (.O (px1901), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[17]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48089z62994.INIT = 32'hD080F0F0;
    LUT5 ix48088z62994 (.O (px1902), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[18]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48088z62994.INIT = 32'hD080F0F0;
    LUT5 ix48087z62994 (.O (px1903), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[19]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48087z62994.INIT = 32'hD080F0F0;
    LUT5 ix48086z62994 (.O (px1904), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[20]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48086z62994.INIT = 32'hD080F0F0;
    LUT5 ix48085z62994 (.O (px1905), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[21]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48085z62994.INIT = 32'hD080F0F0;
    LUT5 ix48084z62994 (.O (px1906), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[22]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48084z62994.INIT = 32'hD080F0F0;
    (* HLUTNM = "LUT62_1_4" *)
    LUT5 ix48083z62994 (.O (px1907), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[23]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48083z62994.INIT = 32'hD080F0F0;
    (* HLUTNM = "LUT62_1_6" *)
    LUT5 ix48082z62994 (.O (px1908), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[24]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48082z62994.INIT = 32'hF2F7F0F0;
    (* HLUTNM = "LUT62_1_30" *)
    LUT5 ix48081z62994 (.O (px1909), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[25]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix48081z62994.INIT = 32'hF2F7F0F0;
    LUT5 ix47093z62994 (.O (px1910), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[26]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix47093z62994.INIT = 32'hF2F7F0F0;
    LUT5 ix47092z62994 (.O (px1911), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[27]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix47092z62994.INIT = 32'hF2F7F0F0;
    LUT5 ix47091z62994 (.O (px1912), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[28]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix47091z62994.INIT = 32'hF2F7F0F0;
    LUT5 ix47090z62994 (.O (px1913), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[29]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix47090z62994.INIT = 32'hF2F7F0F0;
    LUT5 ix47089z62994 (.O (px1914), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[30]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix47089z62994.INIT = 32'hF2F7F0F0;
    LUT5 ix47088z62994 (.O (px1915), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_rec_error_sva[31]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0]), .I4 (
         nx34290z2)) ;
         defparam ix47088z62994.INIT = 32'hF2F7F0F0;
    (* HLUTNM = "LUT62_1_6" *)
    LUT4 ix26190z3404 (.O (nx26190z1), .I0 (nx34290z2), .I1 (\p_fsm_output(10)  
         ), .I2 (main_core_inst_reconstruction_error_rec_error_sva[0]), .I3 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0])) ;
         defparam ix26190z3404.INIT = 16'h082A;
    (* HLUTNM = "LUT62_1_30" *)
    LUT3 ix34290z1354 (.O (nx34290z3), .I0 (\p_fsm_output(10)  ), .I1 (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .I2 (
         main_core_inst_reconstruction_error_for_for_c_mux_nl[0])) ;
         defparam ix34290z1354.INIT = 8'h27;
    (* HLUTNM = "LUT62_1_1" *)
    LUT5 ix38278z2342 (.O (nx38278z1), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (\reconstruction_error_for_acc_3_nl(8)  ), .I3 (
         nx34290z2), .I4 (nx34290z3)) ;
         defparam ix38278z2342.INIT = 32'hAE040404;
    (* HLUTNM = "LUT62_1_1" *)
    LUT5 ix34290z61452 (.O (nx34290z1), .I0 (\fsm_output(9)  ), .I1 (
         \fsm_output(5)  ), .I2 (\reconstruction_error_for_acc_3_nl(8)  ), .I3 (
         nx34290z2), .I4 (nx34290z3)) ;
         defparam ix34290z61452.INIT = 32'h40EAEAEA;
    (* HLUTNM = "LUT62_1_24" *)
    LUT5 ix60483z1314 (.O (nx60483z1), .I0 (nx56495z4), .I1 (p_rst_int), .I2 (
         p_nbus_depth_rsc_addr_1_0[2]), .I3 (nx1399z3), .I4 (\fsm_output(12)  )
         ) ;
         defparam ix60483z1314.INIT = 32'h23100000;
    (* HLUTNM = "LUT62_1_43" *)
    LUT5 ix59486z1314 (.O (nx59486z1), .I0 (\for_1_i_7_0_sva_4(4)  ), .I1 (
         p_nbus_depth_rsc_addr_1_0[2]), .I2 (nx56495z4), .I3 (nx1399z3), .I4 (
         \fsm_output(12)  )) ;
         defparam ix59486z1314.INIT = 32'hA6AA0000;
    DSP48E1 z_out_multu32_0_p_mult0_DSP48E1_0 (.BCOUT ({nx6176z16,nx6176z17,
            nx6176z18,nx6176z19,nx6176z20,nx6176z21,nx6176z22,nx6176z23,
            nx6176z24,nx6176z25,nx6176z26,nx6176z27,nx6176z28,nx6176z29,
            nx6176z30,nx6176z31,nx6176z32,nx6176z33}), .P ({\$dummy [31],
            \$dummy [32],\$dummy [33],\$dummy [34],\$dummy [35],\$dummy [36],
            \$dummy [37],\$dummy [38],\$dummy [39],\$dummy [40],\$dummy [41],
            \$dummy [42],\$dummy [43],\$dummy [44],\$dummy [45],\$dummy [46],
            \$dummy [47],\$dummy [48],\$dummy [49],\$dummy [50],\$dummy [51],
            \$dummy [52],\$dummy [53],\$dummy [54],\$dummy [55],\$dummy [56],
            \$dummy [57],\$dummy [58],\$dummy [59],\$dummy [60],\$dummy [61],
            \z_out(16)  ,\z_out(15)  ,\z_out(14)  ,\z_out(13)  ,\z_out(12)  ,
            \z_out(11)  ,\z_out(10)  ,\z_out(9)  ,\p_z_out(8)  ,\p_z_out(7)  ,
            \p_z_out(6)  ,\p_z_out(5)  ,\p_z_out(4)  ,\p_z_out(3)  ,\p_z_out(2)  
            ,\p_z_out(1)  ,\p_z_out(0)  }), .PCOUT ({nx6176z34,nx6176z35,
            nx6176z36,nx6176z37,nx6176z38,nx6176z39,nx6176z40,nx6176z41,
            nx6176z42,nx6176z43,nx6176z44,nx6176z45,nx6176z46,nx6176z47,
            nx6176z48,nx6176z49,nx6176z50,nx6176z51,nx6176z52,nx6176z53,
            nx6176z54,nx6176z55,nx6176z56,nx6176z57,nx6176z58,nx6176z59,
            nx6176z60,nx6176z61,nx6176z62,nx6176z63,nx6176z64,nx6176z65,
            nx6176z66,nx6176z67,nx6176z68,nx6176z69,nx6176z70,nx6176z71,
            nx6176z72,nx6176z73,nx6176z74,nx6176z75,nx6176z76,nx6176z77,
            nx6176z78,nx6176z79,nx6176z80,nx6176z81}), .A ({px1302,px1302,px1302
            ,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,nx10394z1,nx10394z2,nx10394z3,nx10394z4,nx10394z5,nx10394z6,
            nx10394z7,nx10394z8,nx10394z9,nx10394z11,nx10394z13,nx10394z15,
            nx10394z17,nx10394z19,nx10394z21,nx10394z23,nx10394z25}), .ALUMODE (
            {px1302,px1302,px1302,px1302}), .B ({px1302,nx10394z27,nx10394z28,
            nx10394z29,nx10394z30,nx10394z31,nx10394z32,nx10394z33,nx10394z34,
            nx10394z35,nx10394z36,nx10394z37,nx10394z38,nx10394z39,nx10394z40,
            nx10394z41,nx10394z42,nx10394z43}), .C ({px1302,px1302,px1302,px1302
            ,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302}), .CARRYCASCIN (
            px1302), .CARRYIN (px1302), .CARRYINSEL ({px1302,px1302,px1302}), .CEA1 (
            px1302), .CEA2 (px1302), .CEAD (px1302), .CEALUMODE (px1302), .CEB1 (
            px1302), .CEB2 (px1302), .CEC (px1302), .CECARRYIN (px1302), .CECTRL (
            px1302), .CED (px1302), .CEINMODE (px1302), .CEM (px1302), .CEP (
            px1302), .CLK (px1302), .D ({px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302}), .INMODE ({px1302,px1302,px1302,px1302,px1302}), .MULTSIGNIN (
            px1918), .OPMODE ({px1302,px1302,px1302,px1302,px1918,px1302,px1918}
            ), .RSTA (px1302), .RSTALLCARRYIN (px1302), .RSTALUMODE (px1302), .RSTB (
            px1302), .RSTC (px1302), .RSTCTRL (px1302), .RSTD (px1302), .RSTINMODE (
            px1302), .RSTM (px1302), .RSTP (px1302)) ;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.ACASCREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.ADREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.ALUMODEREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.AREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.AUTORESET_PATDET = "NO_RESET";
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.A_INPUT = "DIRECT";
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.BCASCREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.BREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.B_INPUT = "DIRECT";
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.CARRYINREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.CARRYINSELREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.CREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.DREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.INMODEREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.MREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.OPMODEREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.PREG = 0;
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.SEL_MASK = "MASK";
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.SEL_PATTERN = "PATTERN";
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.USE_DPORT = "FALSE";
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.USE_MULT = "MULTIPLY";
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.USE_PATTERN_DETECT = "NO_PATDET";
            defparam z_out_multu32_0_p_mult0_DSP48E1_0.USE_SIMD = "ONE48";
    DSP48E1 z_out_multu32_0_p_mult1_DSP48E1_1 (.PCOUT ({nx42790z16,nx42790z17,
            nx42790z18,nx42790z19,nx42790z20,nx42790z21,nx42790z22,nx42790z23,
            nx42790z24,nx42790z25,nx42790z26,nx42790z27,nx42790z28,nx42790z29,
            nx42790z30,nx42790z31,nx42790z32,nx42790z33,nx42790z34,nx42790z35,
            nx42790z36,nx42790z37,nx42790z38,nx42790z39,nx42790z40,nx42790z41,
            nx42790z42,nx42790z43,nx42790z44,nx42790z45,nx42790z46,nx42790z47,
            nx42790z48,nx42790z49,nx42790z50,nx42790z51,nx42790z52,nx42790z53,
            nx42790z54,nx42790z55,nx42790z56,nx42790z57,nx42790z58,nx42790z59,
            nx42790z60,nx42790z61,nx42790z62,nx42790z63}), .A ({px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,nx6176z1,nx6176z2,nx6176z3,nx6176z4,
            nx6176z5,nx6176z6,nx6176z7,nx6176z8,nx6176z9,nx6176z10,nx6176z11,
            nx6176z12,nx6176z13,nx6176z14,nx6176z15}), .ALUMODE ({px1302,px1302,
            px1302,px1302}), .BCIN ({nx6176z16,nx6176z17,nx6176z18,nx6176z19,
            nx6176z20,nx6176z21,nx6176z22,nx6176z23,nx6176z24,nx6176z25,
            nx6176z26,nx6176z27,nx6176z28,nx6176z29,nx6176z30,nx6176z31,
            nx6176z32,nx6176z33}), .C ({px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302}), .CARRYCASCIN (
            px1302), .CARRYIN (px1302), .CARRYINSEL ({px1302,px1302,px1302}), .CEA1 (
            px1302), .CEA2 (px1302), .CEAD (px1302), .CEALUMODE (px1302), .CEB1 (
            px1302), .CEB2 (px1302), .CEC (px1302), .CECARRYIN (px1302), .CECTRL (
            px1302), .CED (px1302), .CEINMODE (px1302), .CEM (px1302), .CEP (
            px1302), .CLK (px1302), .D ({px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302}), .INMODE ({px1302,px1302,px1302,px1302,px1302}), .MULTSIGNIN (
            px1918), .OPMODE ({px1918,px1302,px1918,px1302,px1918,px1302,px1918}
            ), .PCIN ({nx6176z34,nx6176z35,nx6176z36,nx6176z37,nx6176z38,
            nx6176z39,nx6176z40,nx6176z41,nx6176z42,nx6176z43,nx6176z44,
            nx6176z45,nx6176z46,nx6176z47,nx6176z48,nx6176z49,nx6176z50,
            nx6176z51,nx6176z52,nx6176z53,nx6176z54,nx6176z55,nx6176z56,
            nx6176z57,nx6176z58,nx6176z59,nx6176z60,nx6176z61,nx6176z62,
            nx6176z63,nx6176z64,nx6176z65,nx6176z66,nx6176z67,nx6176z68,
            nx6176z69,nx6176z70,nx6176z71,nx6176z72,nx6176z73,nx6176z74,
            nx6176z75,nx6176z76,nx6176z77,nx6176z78,nx6176z79,nx6176z80,
            nx6176z81}), .RSTA (px1302), .RSTALLCARRYIN (px1302), .RSTALUMODE (
            px1302), .RSTB (px1302), .RSTC (px1302), .RSTCTRL (px1302), .RSTD (
            px1302), .RSTINMODE (px1302), .RSTM (px1302), .RSTP (px1302)) ;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.ACASCREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.ADREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.ALUMODEREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.AREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.AUTORESET_PATDET = "NO_RESET";
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.A_INPUT = "DIRECT";
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.BCASCREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.BREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.B_INPUT = "CASCADE";
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.CARRYINREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.CARRYINSELREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.CREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.DREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.INMODEREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.MREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.OPMODEREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.PREG = 0;
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.SEL_MASK = "MASK";
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.SEL_PATTERN = "PATTERN";
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.USE_DPORT = "FALSE";
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.USE_MULT = "MULTIPLY";
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.USE_PATTERN_DETECT = "NO_PATDET";
            defparam z_out_multu32_0_p_mult1_DSP48E1_1.USE_SIMD = "ONE48";
    DSP48E1 z_out_multu32_0_p_mult2_DSP48E1_2 (.P ({\$dummy [62],\$dummy [63],
            \$dummy [64],\$dummy [65],\$dummy [66],\$dummy [67],\$dummy [68],
            \$dummy [69],\$dummy [70],\$dummy [71],\$dummy [72],\$dummy [73],
            \$dummy [74],\$dummy [75],\$dummy [76],\$dummy [77],\$dummy [78],
            \$dummy [79],\$dummy [80],\$dummy [81],\$dummy [82],\$dummy [83],
            \$dummy [84],\$dummy [85],\$dummy [86],\$dummy [87],\$dummy [88],
            \$dummy [89],\$dummy [90],\$dummy [91],\$dummy [92],\$dummy [93],
            \$dummy [94],\z_out(31)  ,\z_out(30)  ,\z_out(29)  ,\z_out(28)  ,
            \z_out(27)  ,\z_out(26)  ,\z_out(25)  ,\z_out(24)  ,\z_out(23)  ,
            \z_out(22)  ,\z_out(21)  ,\z_out(20)  ,\z_out(19)  ,\z_out(18)  ,
            main_core_inst_z_out[31]}), .A ({px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,nx10394z1,
            nx10394z2,nx10394z3,nx10394z4,nx10394z5,nx10394z6,nx10394z7,
            nx10394z8,nx10394z9,nx10394z11,nx10394z13,nx10394z15,nx10394z17,
            nx10394z19,nx10394z21,nx10394z23,nx10394z25}), .ALUMODE ({px1302,
            px1302,px1302,px1302}), .B ({px1302,px1302,px1302,nx42790z1,
            nx42790z2,nx42790z3,nx42790z4,nx42790z5,nx42790z6,nx42790z7,
            nx42790z8,nx42790z9,nx42790z10,nx42790z11,nx42790z12,nx42790z13,
            nx42790z14,nx42790z15}), .C ({px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302}), .CARRYCASCIN (
            px1302), .CARRYIN (px1302), .CARRYINSEL ({px1302,px1302,px1302}), .CEA1 (
            px1302), .CEA2 (px1302), .CEAD (px1302), .CEALUMODE (px1302), .CEB1 (
            px1302), .CEB2 (px1302), .CEC (px1302), .CECARRYIN (px1302), .CECTRL (
            px1302), .CED (px1302), .CEINMODE (px1302), .CEM (px1302), .CEP (
            px1302), .CLK (px1302), .D ({px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,px1302,
            px1302,px1302}), .INMODE ({px1302,px1302,px1302,px1302,px1302}), .MULTSIGNIN (
            px1918), .OPMODE ({px1302,px1302,px1918,px1302,px1918,px1302,px1918}
            ), .PCIN ({nx42790z16,nx42790z17,nx42790z18,nx42790z19,nx42790z20,
            nx42790z21,nx42790z22,nx42790z23,nx42790z24,nx42790z25,nx42790z26,
            nx42790z27,nx42790z28,nx42790z29,nx42790z30,nx42790z31,nx42790z32,
            nx42790z33,nx42790z34,nx42790z35,nx42790z36,nx42790z37,nx42790z38,
            nx42790z39,nx42790z40,nx42790z41,nx42790z42,nx42790z43,nx42790z44,
            nx42790z45,nx42790z46,nx42790z47,nx42790z48,nx42790z49,nx42790z50,
            nx42790z51,nx42790z52,nx42790z53,nx42790z54,nx42790z55,nx42790z56,
            nx42790z57,nx42790z58,nx42790z59,nx42790z60,nx42790z61,nx42790z62,
            nx42790z63}), .RSTA (px1302), .RSTALLCARRYIN (px1302), .RSTALUMODE (
            px1302), .RSTB (px1302), .RSTC (px1302), .RSTCTRL (px1302), .RSTD (
            px1302), .RSTINMODE (px1302), .RSTM (px1302), .RSTP (px1302)) ;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.ACASCREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.ADREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.ALUMODEREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.AREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.AUTORESET_PATDET = "NO_RESET";
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.A_INPUT = "DIRECT";
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.BCASCREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.BREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.B_INPUT = "DIRECT";
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.CARRYINREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.CARRYINSELREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.CREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.DREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.INMODEREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.MREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.OPMODEREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.PREG = 0;
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.SEL_MASK = "MASK";
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.SEL_PATTERN = "PATTERN";
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.USE_DPORT = "FALSE";
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.USE_MULT = "MULTIPLY";
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.USE_PATTERN_DETECT = "NO_PATDET";
            defparam z_out_multu32_0_p_mult2_DSP48E1_2.USE_SIMD = "ONE48";
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_0 (.O (nx25626z1), .CI (px1302), .DI (
          nx25625z1), .S (nx25625z2)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_1 (.O (nx25627z1), .CI (nx25626z1)
          , .DI (nx25626z2), .S (nx25626z3)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_2 (.O (nx25628z1), .CI (nx25627z1)
          , .DI (nx25627z2), .S (nx25627z3)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_3 (.O (nx25629z1), .CI (nx25628z1)
          , .DI (nx25628z2), .S (nx25628z3)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_4 (.O (nx25630z1), .CI (nx25629z1)
          , .DI (nx25629z2), .S (nx25629z3)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_5 (.O (nx25631z1), .CI (nx25630z1)
          , .DI (px1302), .S (nx25630z2)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_6 (.O (nx25632z1), .CI (nx25631z1)
          , .DI (px1302), .S (nx25631z2)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_7 (.O (nx25633z1), .CI (nx25632z1)
          , .DI (px1302), .S (nx25632z2)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_8 (.O (nx25634z1), .CI (nx25633z1)
          , .DI (px1302), .S (nx25633z2)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_9 (.O (nx55666z1), .CI (nx25634z1)
          , .DI (px1302), .S (nx25634z2)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_10 (.O (nx55667z1), .CI (nx55666z1
          ), .DI (px1302), .S (nx55666z2)) ;
    MUXCY image_net_rsci_addr_d_add13_4_muxcy_11 (.O (nx40591z1), .CI (nx55667z1
          ), .DI (px1302), .S (nx55667z2)) ;
    MUXCY z_out_2_add8_5_muxcy_0 (.O (nx11511z1), .CI (px1302), .DI (nx11510z2)
          , .S (nx11510z3)) ;
    MUXCY z_out_2_add8_5_muxcy_1 (.O (nx11512z1), .CI (nx11511z1), .DI (
          \p_for_for_mux1h_2_nl(1)  ), .S (nx11511z2)) ;
    MUXCY z_out_2_add8_5_muxcy_2 (.O (nx11513z1), .CI (nx11512z1), .DI (
          nx11512z2), .S (nx11512z3)) ;
    MUXCY z_out_2_add8_5_muxcy_3 (.O (nx11514z1), .CI (nx11513z1), .DI (
          \p_for_for_mux1h_2_nl(1)  ), .S (nx11513z2)) ;
    MUXCY z_out_2_add8_5_muxcy_4 (.O (nx11515z1), .CI (nx11514z1), .DI (
          nx11510z2), .S (nx11514z2)) ;
    MUXCY z_out_2_add8_5_muxcy_5 (.O (nx11516z1), .CI (nx11515z1), .DI (
          nx11510z2), .S (nx11515z2)) ;
    MUXCY z_out_2_add8_5_muxcy_6 (.O (nx48644z1), .CI (nx11516z1), .DI (
          \p_for_for_mux1h_2_nl(1)  ), .S (nx11516z2)) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_0 (.O (nx42708z1), .CI (px1302
          ), .DI (\p_z_out(0)  ), .S (nx42707z1)) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_1 (.O (nx42709z1), .CI (
          nx42708z1), .DI (\p_z_out(1)  ), .S (nx42708z2)) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_2 (.O (nx42710z1), .CI (
          nx42709z1), .DI (\p_z_out(2)  ), .S (nx42709z2)) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_3 (.O (nx42711z1), .CI (
          nx42710z1), .DI (\p_z_out(3)  ), .S (nx42710z2)) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_4 (.O (nx42712z1), .CI (
          nx42711z1), .DI (\p_z_out(4)  ), .S (nx42711z2)) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_5 (.O (nx42713z1), .CI (
          nx42712z1), .DI (px1302), .S (\p_z_out(5)  )) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_6 (.O (nx42714z1), .CI (
          nx42713z1), .DI (px1302), .S (\p_z_out(6)  )) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_7 (.O (nx42715z1), .CI (
          nx42714z1), .DI (px1302), .S (\p_z_out(7)  )) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_8 (.O (nx42716z1), .CI (
          nx42715z1), .DI (px1302), .S (\p_z_out(8)  )) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_9 (.O (nx18476z1), .CI (
          nx42716z1), .DI (px1302), .S (\z_out(9)  )) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_10 (.O (nx18475z1), .CI (
          nx18476z1), .DI (px1302), .S (\z_out(10)  )) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_11 (.O (nx18474z1), .CI (
          nx18475z1), .DI (px1302), .S (\z_out(11)  )) ;
    MUXCY for_for_else_acc_itm_2_add14_14i1_muxcy_12 (.O (nx18473z1), .CI (
          nx18474z1), .DI (px1302), .S (\z_out(12)  )) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_0 (.O (nx12066z1), .CI (
          px1302), .DI (nx12067z1), .S (nx12067z2)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_1 (.O (nx12065z1), .CI (
          nx12066z1), .DI (nx12066z2), .S (nx12066z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_2 (.O (nx12064z1), .CI (
          nx12065z1), .DI (nx12065z2), .S (nx12065z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_3 (.O (nx12063z1), .CI (
          nx12064z1), .DI (nx12064z2), .S (nx12064z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_4 (.O (nx12062z1), .CI (
          nx12063z1), .DI (nx12063z2), .S (nx12063z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_5 (.O (nx12061z1), .CI (
          nx12062z1), .DI (nx12062z2), .S (nx12062z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_6 (.O (nx12060z1), .CI (
          nx12061z1), .DI (nx12061z2), .S (nx12061z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_7 (.O (nx12059z1), .CI (
          nx12060z1), .DI (nx12060z2), .S (nx12060z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_8 (.O (nx12058z1), .CI (
          nx12059z1), .DI (nx12059z2), .S (nx12059z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_9 (.O (nx36666z1), .CI (
          nx12058z1), .DI (nx12058z2), .S (nx12058z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_10 (.O (nx36665z1), .CI (
          nx36666z1), .DI (nx36666z2), .S (nx36666z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_11 (.O (nx36664z1), .CI (
          nx36665z1), .DI (nx36665z2), .S (nx36665z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_12 (.O (nx36663z1), .CI (
          nx36664z1), .DI (nx36664z2), .S (nx36664z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_13 (.O (nx36662z1), .CI (
          nx36663z1), .DI (nx36663z2), .S (nx36663z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_14 (.O (nx36661z1), .CI (
          nx36662z1), .DI (nx36662z2), .S (nx36662z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_15 (.O (nx36660z1), .CI (
          nx36661z1), .DI (nx36661z2), .S (nx36661z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_16 (.O (nx36659z1), .CI (
          nx36660z1), .DI (nx36660z2), .S (nx36660z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_17 (.O (nx36658z1), .CI (
          nx36659z1), .DI (nx36659z2), .S (nx36659z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_18 (.O (nx36657z1), .CI (
          nx36658z1), .DI (nx36658z2), .S (nx36658z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_19 (.O (nx35669z1), .CI (
          nx36657z1), .DI (nx36657z2), .S (nx36657z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_20 (.O (nx35668z1), .CI (
          nx35669z1), .DI (nx35669z2), .S (nx35669z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_21 (.O (nx35667z1), .CI (
          nx35668z1), .DI (nx35668z2), .S (nx35668z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_22 (.O (nx35666z1), .CI (
          nx35667z1), .DI (nx35667z2), .S (nx35667z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_23 (.O (nx35665z1), .CI (
          nx35666z1), .DI (nx35666z2), .S (nx35666z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_24 (.O (nx35664z1), .CI (
          nx35665z1), .DI (nx35665z2), .S (nx35665z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_25 (.O (nx35663z1), .CI (
          nx35664z1), .DI (nx35664z2), .S (nx35664z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_26 (.O (nx35662z1), .CI (
          nx35663z1), .DI (nx35663z2), .S (nx35663z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_27 (.O (nx35661z1), .CI (
          nx35662z1), .DI (nx35662z2), .S (nx35662z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_28 (.O (nx35660z1), .CI (
          nx35661z1), .DI (nx35661z2), .S (nx35661z3)) ;
    MUXCY reconstruction_error_for_acc_nl_add31_11_muxcy_29 (.O (nx34672z1), .CI (
          nx35660z1), .DI (nx35660z2), .S (nx35660z3)) ;
    MUXCY muxcy_0_3 (.O (nx39520z1), .CI (nx39519z1), .DI (nx39519z2), .S (
          nx39519z1)) ;
    MUXCY muxcy_0_4 (.O (nx39521z1), .CI (nx39520z1), .DI (nx39520z2), .S (
          nx39520z3)) ;
    MUXCY muxcy_0_5 (.O (nx39522z1), .CI (nx39521z1), .DI (nx39521z2), .S (
          nx39521z3)) ;
    MUXCY muxcy_0_6 (.O (nx39523z1), .CI (nx39522z1), .DI (nx39522z2), .S (
          nx39522z3)) ;
    MUXCY muxcy_0_7 (.O (nx39524z1), .CI (nx39523z1), .DI (nx39523z2), .S (
          nx39523z3)) ;
    MUXCY muxcy_0_8 (.O (nx50036z1), .CI (nx39524z1), .DI (nx39524z2), .S (
          nx39524z3)) ;
    MUXCY z_out_6_add33_6_muxcy_0 (.O (nx42643z1), .CI (not_fsm_output_8), .DI (
          nx17517z1), .S (nx42644z1)) ;
    MUXCY z_out_6_add33_6_muxcy_1 (.O (nx42642z1), .CI (nx42643z1), .DI (
          nx17518z1), .S (nx42643z2)) ;
    MUXCY z_out_6_add33_6_muxcy_2 (.O (nx42641z1), .CI (nx42642z1), .DI (
          nx17519z1), .S (nx42642z2)) ;
    MUXCY z_out_6_add33_6_muxcy_3 (.O (nx42640z1), .CI (nx42641z1), .DI (
          nx17520z1), .S (nx42641z2)) ;
    MUXCY z_out_6_add33_6_muxcy_4 (.O (nx42639z1), .CI (nx42640z1), .DI (
          nx17521z1), .S (nx42640z2)) ;
    MUXCY z_out_6_add33_6_muxcy_5 (.O (nx42638z1), .CI (nx42639z1), .DI (
          nx17522z1), .S (nx42639z2)) ;
    MUXCY z_out_6_add33_6_muxcy_6 (.O (nx42637z1), .CI (nx42638z1), .DI (
          nx17523z1), .S (nx42638z2)) ;
    MUXCY z_out_6_add33_6_muxcy_7 (.O (nx42636z1), .CI (nx42637z1), .DI (
          nx17524z1), .S (nx42637z2)) ;
    MUXCY z_out_6_add33_6_muxcy_8 (.O (nx42635z1), .CI (nx42636z1), .DI (
          nx17525z1), .S (nx42636z2)) ;
    MUXCY z_out_6_add33_6_muxcy_9 (.O (nx47695z1), .CI (nx42635z1), .DI (
          nx17526z1), .S (nx42635z2)) ;
    MUXCY z_out_6_add33_6_muxcy_10 (.O (nx47694z1), .CI (nx47695z1), .DI (
          nx32918z1), .S (nx47695z2)) ;
    MUXCY z_out_6_add33_6_muxcy_11 (.O (nx47693z1), .CI (nx47694z1), .DI (
          nx32919z1), .S (nx47694z2)) ;
    MUXCY z_out_6_add33_6_muxcy_12 (.O (nx47692z1), .CI (nx47693z1), .DI (
          nx32920z1), .S (nx47693z2)) ;
    MUXCY z_out_6_add33_6_muxcy_13 (.O (nx47691z1), .CI (nx47692z1), .DI (
          nx32921z1), .S (nx47692z2)) ;
    MUXCY z_out_6_add33_6_muxcy_14 (.O (nx47690z1), .CI (nx47691z1), .DI (
          nx32922z1), .S (nx47691z2)) ;
    MUXCY z_out_6_add33_6_muxcy_15 (.O (nx47689z1), .CI (nx47690z1), .DI (
          nx32923z1), .S (nx47690z2)) ;
    MUXCY z_out_6_add33_6_muxcy_16 (.O (nx47688z1), .CI (nx47689z1), .DI (
          nx32924z1), .S (nx47689z2)) ;
    MUXCY z_out_6_add33_6_muxcy_17 (.O (nx47687z1), .CI (nx47688z1), .DI (
          nx32925z1), .S (nx47688z2)) ;
    MUXCY z_out_6_add33_6_muxcy_18 (.O (nx47686z1), .CI (nx47687z1), .DI (
          nx32926z1), .S (nx47687z2)) ;
    MUXCY z_out_6_add33_6_muxcy_19 (.O (nx46698z1), .CI (nx47686z1), .DI (
          nx32927z1), .S (nx47686z2)) ;
    MUXCY z_out_6_add33_6_muxcy_20 (.O (nx46697z1), .CI (nx46698z1), .DI (
          nx33915z1), .S (nx46698z2)) ;
    MUXCY z_out_6_add33_6_muxcy_21 (.O (nx46696z1), .CI (nx46697z1), .DI (
          nx33916z1), .S (nx46697z2)) ;
    MUXCY z_out_6_add33_6_muxcy_22 (.O (nx46695z1), .CI (nx46696z1), .DI (
          nx33917z1), .S (nx46696z2)) ;
    MUXCY z_out_6_add33_6_muxcy_23 (.O (nx46694z1), .CI (nx46695z1), .DI (
          nx33918z1), .S (nx46695z2)) ;
    MUXCY z_out_6_add33_6_muxcy_24 (.O (nx46693z1), .CI (nx46694z1), .DI (
          nx33919z1), .S (nx46694z2)) ;
    MUXCY z_out_6_add33_6_muxcy_25 (.O (nx46692z1), .CI (nx46693z1), .DI (
          nx33920z1), .S (nx46693z2)) ;
    MUXCY z_out_6_add33_6_muxcy_26 (.O (nx46691z1), .CI (nx46692z1), .DI (
          nx33921z1), .S (nx46692z2)) ;
    MUXCY z_out_6_add33_6_muxcy_27 (.O (nx46690z1), .CI (nx46691z1), .DI (
          nx33922z1), .S (nx46691z2)) ;
    MUXCY z_out_6_add33_6_muxcy_28 (.O (nx46689z1), .CI (nx46690z1), .DI (
          nx33923z1), .S (nx46690z2)) ;
    MUXCY z_out_6_add33_6_muxcy_29 (.O (nx45701z1), .CI (nx46689z1), .DI (
          nx33924z1), .S (nx46689z2)) ;
    MUXCY z_out_6_add33_6_muxcy_30 (.O (nx45700z1), .CI (nx45701z1), .DI (
          nx34912z1), .S (nx45701z2)) ;
    MUXCY reconstruction_error_for_acc_3_nl_add9_1_muxcy_0 (.O (nx7972z1), .CI (
          \reconstruction_error_for_acc_3_nl_0n0s2(0)  ), .DI (nx7971z1), .S (
          p_nbus_depth_rsc_addr_1_0[0])) ;
    MUXCY reconstruction_error_for_acc_3_nl_add9_1_muxcy_1 (.O (nx7973z1), .CI (
          nx7972z1), .DI (nx7972z2), .S (nx7972z3)) ;
    MUXCY reconstruction_error_for_acc_3_nl_add9_1_muxcy_2 (.O (nx7974z1), .CI (
          nx7973z1), .DI (nx7973z2), .S (nx7973z4)) ;
    MUXCY reconstruction_error_for_acc_3_nl_add9_1_muxcy_3 (.O (nx7975z1), .CI (
          nx7974z1), .DI (nx7974z2), .S (nx7974z4)) ;
    MUXCY reconstruction_error_for_acc_3_nl_add9_1_muxcy_4 (.O (nx7976z1), .CI (
          nx7975z1), .DI (nx7975z2), .S (nx7975z5)) ;
    MUXCY reconstruction_error_for_acc_3_nl_add9_1_muxcy_5 (.O (nx7977z1), .CI (
          nx7976z1), .DI (nx7976z2), .S (nx7976z6)) ;
    MUXCY reconstruction_error_for_acc_3_nl_add9_1_muxcy_6 (.O (nx52183z1), .CI (
          nx7977z1), .DI (nx7977z2), .S (nx7977z6)) ;
    MUXCY modgen_add_4_muxcy_0 (.O (nx33895z1), .CI (px1302), .DI (px1658), .S (
          nx33896z1)) ;
    MUXCY modgen_add_4_muxcy_1 (.O (nx33894z1), .CI (nx33895z1), .DI (px1656), .S (
          nx33895z2)) ;
    MUXCY modgen_add_4_muxcy_2 (.O (nx33893z1), .CI (nx33894z1), .DI (px1654), .S (
          nx33894z2)) ;
    MUXCY modgen_add_4_muxcy_3 (.O (nx33892z1), .CI (nx33893z1), .DI (px1652), .S (
          nx33893z2)) ;
    MUXCY modgen_add_4_muxcy_4 (.O (nx33891z1), .CI (nx33892z1), .DI (px1650), .S (
          nx33892z2)) ;
    MUXCY modgen_add_4_muxcy_5 (.O (nx33890z1), .CI (nx33891z1), .DI (px1648), .S (
          nx33891z2)) ;
    MUXCY modgen_add_4_muxcy_6 (.O (nx33889z1), .CI (nx33890z1), .DI (px1646), .S (
          nx33890z2)) ;
    MUXCY modgen_add_4_muxcy_7 (.O (nx33888z1), .CI (nx33889z1), .DI (px1644), .S (
          nx33889z2)) ;
    MUXCY modgen_add_4_muxcy_8 (.O (nx33887z1), .CI (nx33888z1), .DI (px1642), .S (
          nx33888z2)) ;
    MUXCY modgen_add_4_muxcy_9 (.O (nx23309z1), .CI (nx33887z1), .DI (nx26274z1)
          , .S (nx33887z2)) ;
    MUXCY modgen_add_4_muxcy_10 (.O (nx23310z1), .CI (nx23309z1), .DI (nx38386z1
          ), .S (nx23309z2)) ;
    MUXCY modgen_add_4_muxcy_11 (.O (nx23311z1), .CI (nx23310z1), .DI (nx38387z1
          ), .S (nx23310z2)) ;
    MUXCY modgen_add_4_muxcy_12 (.O (nx23312z1), .CI (nx23311z1), .DI (nx38388z1
          ), .S (nx23311z2)) ;
    MUXCY ix456_muxcy_0 (.O (nx42832z1), .CI (px1302), .DI (
          main_core_inst_for_for_j_8_0_sva_3[0]), .S (nx42831z1)) ;
    MUXCY ix456_muxcy_1 (.O (nx42833z1), .CI (nx42832z1), .DI (
          main_core_inst_for_for_j_8_0_sva_3[1]), .S (nx42832z2)) ;
    MUXCY ix456_muxcy_2 (.O (nx42834z1), .CI (nx42833z1), .DI (
          main_core_inst_for_for_j_8_0_sva_3[2]), .S (nx42833z2)) ;
    MUXCY ix456_muxcy_3 (.O (nx42835z1), .CI (nx42834z1), .DI (
          main_core_inst_for_for_j_8_0_sva_3[3]), .S (nx42834z2)) ;
    MUXCY ix456_muxcy_4 (.O (nx42836z1), .CI (nx42835z1), .DI (
          main_core_inst_for_for_j_8_0_sva_3[4]), .S (nx42835z2)) ;
    MUXCY ix456_muxcy_5 (.O (nx42837z1), .CI (nx42836z1), .DI (
          main_core_inst_for_for_j_8_0_sva_3[5]), .S (nx42836z2)) ;
    MUXCY ix456_muxcy_6 (.O (nx42838z1), .CI (nx42837z1), .DI (
          main_core_inst_for_for_j_8_0_sva_3[6]), .S (nx42837z2)) ;
    MUXCY ix456_muxcy_7 (.O (nx42839z1), .CI (nx42838z1), .DI (px1302), .S (
          main_core_inst_for_for_j_8_0_sva_3[5])) ;
    MUXCY ix486_muxcy_0 (.O (nx60385z1), .CI (px1302), .DI (\a(0)  ), .S (
          nx60386z1)) ;
    MUXCY ix486_muxcy_1 (.O (nx60384z1), .CI (nx60385z1), .DI (\a(1)  ), .S (
          nx60385z2)) ;
    MUXCY ix486_muxcy_2 (.O (nx60383z1), .CI (nx60384z1), .DI (\a(2)  ), .S (
          nx60384z2)) ;
    MUXCY ix486_muxcy_3 (.O (nx60382z1), .CI (nx60383z1), .DI (\a(3)  ), .S (
          nx60383z2)) ;
    MUXCY ix486_muxcy_4 (.O (nx60381z1), .CI (nx60382z1), .DI (\a(4)  ), .S (
          nx60382z2)) ;
    MUXCY ix486_muxcy_5 (.O (nx60380z1), .CI (nx60381z1), .DI (\a(5)  ), .S (
          nx60381z2)) ;
    MUXCY ix486_muxcy_6 (.O (nx60379z1), .CI (nx60380z1), .DI (\a(6)  ), .S (
          nx60380z2)) ;
    MUXCY ix486_muxcy_7 (.O (nx60378z1), .CI (nx60379z1), .DI (\a(7)  ), .S (
          nx60379z2)) ;
    MUXCY ix486_muxcy_8 (.O (nx60377z1), .CI (nx60378z1), .DI (\a(8)  ), .S (
          nx60378z2)) ;
    MUXCY ix486_muxcy_9 (.O (nx41749z1), .CI (nx60377z1), .DI (\a(9)  ), .S (
          nx60377z2)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(8)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[0]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx21850z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(7)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[1]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx22847z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(6)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[2]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx23844z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(5)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[3]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx24841z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(4)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[4]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx25838z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(3)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[5]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx26835z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(2)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[6]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx27832z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(1)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[7]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx57639z1), .R (p_rst_int)) ;
    FDRE \reg_for_1_for_j_8_0_sva_4(0)  (.Q (
         main_core_inst_for_1_for_j_8_0_sva_4[8]), .C (p_clk_int), .CE (
         nx39519z3), .D (nx56642z1), .R (p_rst_int)) ;
    FDRE reg_for_1_for_slc_for_1_for_acc_7_itm_1 (.Q (
         for_1_for_slc_for_1_for_acc_7_itm_1), .C (p_clk_int), .CE (nx39519z3), 
         .D (main_core_inst_z_out_2[7]), .R (p_rst_int)) ;
    FDRE reg_exit_reconstruction_error_for_for_sva_1 (.Q (
         exit_reconstruction_error_for_for_sva_1), .C (p_clk_int), .CE (
         nx39519z3), .D (nx26190z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(31)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[0]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx4228z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(30)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[1]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx3231z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(29)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[2]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx1235z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(28)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[3]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx238z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(27)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[4]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx64777z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(26)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[5]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx63780z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(25)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[6]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx62783z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(24)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[7]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx61786z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(23)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[8]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx60789z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(22)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[9]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx59792z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(21)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[10]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx58795z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(20)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[11]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx57798z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(19)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[12]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx55802z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(18)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[13]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx54805z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(17)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[14]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx53808z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(16)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[15]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx52811z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(15)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[16]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx51814z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(14)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[17]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx50817z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(13)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[18]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx49820z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(12)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[19]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx48823z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(11)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[20]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx47826z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(10)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[21]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx46829z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(9)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[22]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx5781z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(8)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[23]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx4784z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(7)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[24]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx3787z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(6)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[25]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx2790z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(5)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[26]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx1793z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(4)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[27]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx796z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(3)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[28]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx65335z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(2)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[29]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx64338z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(1)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[30]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx63341z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_lpi_6(0)  (.Q (
         main_core_inst_reconstruction_error_rec_error_lpi_6[31]), .C (p_clk_int
         ), .CE (nx39519z3), .D (nx62344z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(31)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[0]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx29656z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(30)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[1]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx30653z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(29)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[2]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx32649z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(28)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[3]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx33646z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(27)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[4]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx34643z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(26)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[5]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx35640z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(25)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[6]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx36637z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(24)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[7]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx37634z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(23)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[8]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx38631z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(22)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[9]), .C (p_clk_int), 
         .CE (nx39519z3), .D (nx39628z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(21)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[10]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx40625z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(20)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[11]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx41622z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(19)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[12]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx43618z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(18)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[13]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx44615z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(17)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[14]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx45612z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(16)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[15]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx46609z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(15)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[16]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx47606z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(14)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[17]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx48603z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(13)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[18]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx49600z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(12)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[19]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx50597z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(11)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[20]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx51594z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(10)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[21]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx52591z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(9)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[22]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx52887z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(8)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[23]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx53884z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(7)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[24]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx54881z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(6)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[25]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx55878z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(5)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[26]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx56875z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(4)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[27]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx57872z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(3)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[28]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx58869z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(2)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[29]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx59866z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(1)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[30]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx60863z1), .R (p_rst_int)) ;
    FDRE \reg_reconstruction_error_rec_error_sva(0)  (.Q (
         main_core_inst_reconstruction_error_rec_error_sva[31]), .C (p_clk_int)
         , .CE (nx39519z3), .D (nx61860z1), .R (p_rst_int)) ;
    FDRE reg_for_for_if_for_for_if_and_itm_1 (.Q (
         for_for_if_for_for_if_and_itm_1), .C (p_clk_int), .CE (nx39519z3), .D (
         nx6053z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(13)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[0]), .C (p_clk_int), .CE (
         nx39519z3), .D (\for_for_else_acc_itm_2_14n1s1(13)  ), .R (p_rst_int)
         ) ;
    FDRE \reg_for_for_else_acc_itm_2(12)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[1]), .C (p_clk_int), .CE (
         nx39519z3), .D (\for_for_else_acc_itm_2_14n1s1(12)  ), .R (p_rst_int)
         ) ;
    FDRE \reg_for_for_else_acc_itm_2(11)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[2]), .C (p_clk_int), .CE (
         nx39519z3), .D (\for_for_else_acc_itm_2_14n1s1(11)  ), .R (p_rst_int)
         ) ;
    FDRE \reg_for_for_else_acc_itm_2(10)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[3]), .C (p_clk_int), .CE (
         nx39519z3), .D (\for_for_else_acc_itm_2_14n1s1(10)  ), .R (p_rst_int)
         ) ;
    FDRE \reg_for_for_else_acc_itm_2(9)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[4]), .C (p_clk_int), .CE (
         nx39519z3), .D (\for_for_else_acc_itm_2_14n1s1(9)  ), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(8)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[5]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[8]), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(7)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[6]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[7]), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(6)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[7]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[6]), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(5)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[8]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[5]), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(4)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[9]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[4]), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(3)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[10]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[3]), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(2)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[11]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[2]), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(1)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[12]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[1]), .R (p_rst_int)) ;
    FDRE \reg_for_for_else_acc_itm_2(0)  (.Q (
         main_core_inst_for_for_else_acc_itm_2[13]), .C (p_clk_int), .CE (
         nx39519z3), .D (main_core_inst_for_for_if_acc_nl[0]), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(8)  (.Q (main_core_inst_for_for_j_8_0_sva_3[6]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx7501z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(7)  (.Q (main_core_inst_for_for_j_8_0_sva_3[5]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx6504z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(6)  (.Q (main_core_inst_for_for_j_8_0_sva_3[4]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx5507z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(5)  (.Q (main_core_inst_for_for_j_8_0_sva_3[3]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx4510z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(4)  (.Q (main_core_inst_for_for_j_8_0_sva_3[2]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx3513z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(3)  (.Q (main_core_inst_for_for_j_8_0_sva_3[1]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx2516z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(2)  (.Q (main_core_inst_for_for_j_8_0_sva_3[0]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx1519z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(1)  (.Q (main_core_inst_for_for_j_8_0_sva_3[7]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx522z1), .R (p_rst_int)) ;
    FDRE \reg_for_for_j_8_0_sva_3(0)  (.Q (main_core_inst_for_for_j_8_0_sva_3[8]
         ), .C (p_clk_int), .CE (nx39519z3), .D (nx65061z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(12)  (.Q (
         p_image_net_rsc_triosy_lz_1_0), .C (p_clk_int), .CE (nx39519z3), .D (
         nx8012z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(11)  (.Q (\fsm_output(12)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (nx7015z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(10)  (.Q (\fsm_output(11)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (\p_fsm_output(10)  ), .R (p_rst_int)
         ) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(9)  (.Q (\p_fsm_output(10)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (nx38278z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(8)  (.Q (\fsm_output(9)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (nx37281z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(7)  (.Q (\fsm_output(8)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (\p_for_for_mux1h_2_nl(1)  ), .R (
         p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(6)  (.Q (
         \p_for_for_mux1h_2_nl(1)  ), .C (p_clk_int), .CE (nx39519z3), .D (
         nx35287z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(5)  (.Q (\fsm_output(6)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (nx34290z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(4)  (.Q (\fsm_output(5)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (nx33293z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(3)  (.Q (\fsm_output(4)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (nx32296z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(2)  (.Q (
         \main_core_core_fsm_inst_fsm_output(3)  ), .C (p_clk_int), .CE (
         nx39519z3), .D (nx31299z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(0)  (.Q (\fsm_output(1)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (nx29305z1), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(1)  (.Q (nx31299z1), .C (
         p_clk_int), .CE (nx39519z3), .D (\fsm_output(1)  ), .R (p_rst_int)) ;
    FDRE \main_core_core_fsm_inst_reg_state_var(13)  (.Q (\fsm_output(0)  ), .C (
         p_clk_int), .CE (nx39519z3), .D (nx9009z1), .R (nx39519z1)) ;
    FDRE \reg_for_1_i_7_0_sva_4(7)  (.Q (nx63944z3), .C (p_clk_int), .CE (
         nx56495z1), .D (nx56495z2), .R (nx39519z1)) ;
    FDRE \reg_for_1_i_7_0_sva_4(6)  (.Q (nx56495z7), .C (p_clk_int), .CE (
         nx56495z1), .D (nx57492z1), .R (nx39519z1)) ;
    FDRE \reg_for_1_i_7_0_sva_4(5)  (.Q (nx64941z4), .C (p_clk_int), .CE (
         nx56495z1), .D (nx58489z1), .R (nx39519z1)) ;
    FDRE \reg_for_1_i_7_0_sva_4(3)  (.Q (nx1399z3), .C (p_clk_int), .CE (
         nx56495z1), .D (nx60483z1), .R (nx39519z1)) ;
    FDRE \reg_for_1_i_7_0_sva_4(2)  (.Q (p_nbus_depth_rsc_addr_1_0[2]), .C (
         p_clk_int), .CE (nx56495z1), .D (nx61480z1), .R (nx39519z1)) ;
endmodule


module inc_32_0 ( cin, a, d, cout, 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(21)  , 
                  \p_for_for_mux1h_2_nl(1)  , 
                  \p_reconstruction_error_for_l_sva_3(30)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(20)  , 
                  \p_reconstruction_error_for_l_sva_3(29)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(19)  , 
                  \p_reconstruction_error_for_l_sva_3(28)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(18)  , 
                  \p_reconstruction_error_for_l_sva_3(27)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(17)  , 
                  \p_reconstruction_error_for_l_sva_3(26)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(16)  , 
                  \p_reconstruction_error_for_l_sva_3(25)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(15)  , 
                  \p_reconstruction_error_for_l_sva_3(24)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(14)  , 
                  \p_reconstruction_error_for_l_sva_3(23)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(13)  , 
                  \p_reconstruction_error_for_l_sva_3(22)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(12)  , 
                  \p_reconstruction_error_for_l_sva_3(21)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(11)  , 
                  \p_reconstruction_error_for_l_sva_3(20)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(10)  , 
                  \p_reconstruction_error_for_l_sva_3(19)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(9)  , 
                  \p_reconstruction_error_for_l_sva_3(18)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(8)  , 
                  \p_reconstruction_error_for_l_sva_3(17)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(7)  , 
                  \p_reconstruction_error_for_l_sva_3(16)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(6)  , 
                  \p_reconstruction_error_for_l_sva_3(15)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(5)  , 
                  \p_reconstruction_error_for_l_sva_3(14)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(4)  , 
                  \p_reconstruction_error_for_l_sva_3(13)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(3)  , 
                  \p_reconstruction_error_for_l_sva_3(12)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(2)  , 
                  \p_reconstruction_error_for_l_sva_3(11)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(1)  , 
                  \p_reconstruction_error_for_l_sva_3(10)  , 
                  \p_reconstruction_error_for_for_c_sva_31_9_2(0)  , 
                  \p_reconstruction_error_for_l_sva_3(9)  , 
                  \p_reconstruction_error_for_l_sva_3(8)  , px2488, 
                  \p_reconstruction_error_for_l_sva_3(7)  , px2489, 
                  \p_reconstruction_error_for_l_sva_3(6)  , px2490, 
                  \p_reconstruction_error_for_l_sva_3(5)  , px2491, 
                  \p_reconstruction_error_for_l_sva_3(4)  , px2492, 
                  \p_reconstruction_error_for_l_sva_3(3)  , px2493, 
                  \p_reconstruction_error_for_l_sva_3(2)  , px2494, 
                  \p_reconstruction_error_for_l_sva_3(1)  , px2495, 
                  \p_reconstruction_error_for_l_sva_3(0)  , px2496 ) ;

    input cin ;
    input [31:0]a ;
    output [31:0]d ;
    output cout ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(21)   ;
    input \p_for_for_mux1h_2_nl(1)   ;
    input \p_reconstruction_error_for_l_sva_3(30)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(20)   ;
    input \p_reconstruction_error_for_l_sva_3(29)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(19)   ;
    input \p_reconstruction_error_for_l_sva_3(28)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(18)   ;
    input \p_reconstruction_error_for_l_sva_3(27)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(17)   ;
    input \p_reconstruction_error_for_l_sva_3(26)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(16)   ;
    input \p_reconstruction_error_for_l_sva_3(25)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(15)   ;
    input \p_reconstruction_error_for_l_sva_3(24)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(14)   ;
    input \p_reconstruction_error_for_l_sva_3(23)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(13)   ;
    input \p_reconstruction_error_for_l_sva_3(22)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(12)   ;
    input \p_reconstruction_error_for_l_sva_3(21)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(11)   ;
    input \p_reconstruction_error_for_l_sva_3(20)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(10)   ;
    input \p_reconstruction_error_for_l_sva_3(19)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(9)   ;
    input \p_reconstruction_error_for_l_sva_3(18)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(8)   ;
    input \p_reconstruction_error_for_l_sva_3(17)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(7)   ;
    input \p_reconstruction_error_for_l_sva_3(16)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(6)   ;
    input \p_reconstruction_error_for_l_sva_3(15)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(5)   ;
    input \p_reconstruction_error_for_l_sva_3(14)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(4)   ;
    input \p_reconstruction_error_for_l_sva_3(13)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(3)   ;
    input \p_reconstruction_error_for_l_sva_3(12)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(2)   ;
    input \p_reconstruction_error_for_l_sva_3(11)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(1)   ;
    input \p_reconstruction_error_for_l_sva_3(10)   ;
    input \p_reconstruction_error_for_for_c_sva_31_9_2(0)   ;
    input \p_reconstruction_error_for_l_sva_3(9)   ;
    input \p_reconstruction_error_for_l_sva_3(8)   ;
    input px2488 ;
    input \p_reconstruction_error_for_l_sva_3(7)   ;
    input px2489 ;
    input \p_reconstruction_error_for_l_sva_3(6)   ;
    input px2490 ;
    input \p_reconstruction_error_for_l_sva_3(5)   ;
    input px2491 ;
    input \p_reconstruction_error_for_l_sva_3(4)   ;
    input px2492 ;
    input \p_reconstruction_error_for_l_sva_3(3)   ;
    input px2493 ;
    input \p_reconstruction_error_for_l_sva_3(2)   ;
    input px2494 ;
    input \p_reconstruction_error_for_l_sva_3(1)   ;
    input px2495 ;
    input \p_reconstruction_error_for_l_sva_3(0)   ;
    input px2496 ;

    wire nx8473z2, nx8473z1, nx8473z3, nx8474z1, nx8474z2, nx8475z1, nx8475z2, 
         nx8476z1, nx8476z2, nx8477z1, nx8477z2, nx8478z1, nx8478z2, nx8479z1, 
         nx8479z2, nx8480z1, nx8480z2, nx8481z1, nx8481z2, nx8482z1, nx8482z2, 
         nx60018z1, nx60018z2, nx60019z1, nx60019z2, nx60020z1, nx60020z2, 
         nx60021z1, nx60021z2, nx60022z1, nx60022z2, nx60023z1, nx60023z2, 
         nx60024z1, nx60024z2, nx60025z1, nx60025z2, nx60026z1, nx60026z2, 
         nx60027z1, nx60027z2, nx61015z1, nx61015z2, nx61016z1, nx61016z2, 
         nx61017z1, nx61017z2, nx61018z1, nx61018z2, nx61019z1, nx61019z2, 
         nx61020z1, nx61020z2, nx61021z1, nx61021z2, nx61022z1, nx61022z2, 
         nx61023z1, nx61023z2, nx61024z1, nx61024z2, nx62012z1, nx62012z2, 
         nx18600z1;



    GND ps_gnd (.G (nx8473z2)) ;
    VCC ps_vcc (.P (nx8473z1)) ;
    XORCY xorcy_0 (.O (d[0]), .CI (nx8473z1), .LI (nx8473z3)) ;
    XORCY xorcy_1 (.O (d[1]), .CI (nx8474z1), .LI (nx8474z2)) ;
    XORCY xorcy_2 (.O (d[2]), .CI (nx8475z1), .LI (nx8475z2)) ;
    XORCY xorcy_3 (.O (d[3]), .CI (nx8476z1), .LI (nx8476z2)) ;
    XORCY xorcy_4 (.O (d[4]), .CI (nx8477z1), .LI (nx8477z2)) ;
    XORCY xorcy_5 (.O (d[5]), .CI (nx8478z1), .LI (nx8478z2)) ;
    XORCY xorcy_6 (.O (d[6]), .CI (nx8479z1), .LI (nx8479z2)) ;
    XORCY xorcy_7 (.O (d[7]), .CI (nx8480z1), .LI (nx8480z2)) ;
    XORCY xorcy_8 (.O (d[8]), .CI (nx8481z1), .LI (nx8481z2)) ;
    XORCY xorcy_9 (.O (d[9]), .CI (nx8482z1), .LI (nx8482z2)) ;
    XORCY xorcy_10 (.O (d[10]), .CI (nx60018z1), .LI (nx60018z2)) ;
    XORCY xorcy_11 (.O (d[11]), .CI (nx60019z1), .LI (nx60019z2)) ;
    XORCY xorcy_12 (.O (d[12]), .CI (nx60020z1), .LI (nx60020z2)) ;
    XORCY xorcy_13 (.O (d[13]), .CI (nx60021z1), .LI (nx60021z2)) ;
    XORCY xorcy_14 (.O (d[14]), .CI (nx60022z1), .LI (nx60022z2)) ;
    XORCY xorcy_15 (.O (d[15]), .CI (nx60023z1), .LI (nx60023z2)) ;
    XORCY xorcy_16 (.O (d[16]), .CI (nx60024z1), .LI (nx60024z2)) ;
    XORCY xorcy_17 (.O (d[17]), .CI (nx60025z1), .LI (nx60025z2)) ;
    XORCY xorcy_18 (.O (d[18]), .CI (nx60026z1), .LI (nx60026z2)) ;
    XORCY xorcy_19 (.O (d[19]), .CI (nx60027z1), .LI (nx60027z2)) ;
    XORCY xorcy_20 (.O (d[20]), .CI (nx61015z1), .LI (nx61015z2)) ;
    XORCY xorcy_21 (.O (d[21]), .CI (nx61016z1), .LI (nx61016z2)) ;
    XORCY xorcy_22 (.O (d[22]), .CI (nx61017z1), .LI (nx61017z2)) ;
    XORCY xorcy_23 (.O (d[23]), .CI (nx61018z1), .LI (nx61018z2)) ;
    XORCY xorcy_24 (.O (d[24]), .CI (nx61019z1), .LI (nx61019z2)) ;
    XORCY xorcy_25 (.O (d[25]), .CI (nx61020z1), .LI (nx61020z2)) ;
    XORCY xorcy_26 (.O (d[26]), .CI (nx61021z1), .LI (nx61021z2)) ;
    XORCY xorcy_27 (.O (d[27]), .CI (nx61022z1), .LI (nx61022z2)) ;
    XORCY xorcy_28 (.O (d[28]), .CI (nx61023z1), .LI (nx61023z2)) ;
    XORCY xorcy_29 (.O (d[29]), .CI (nx61024z1), .LI (nx61024z2)) ;
    XORCY xorcy_30 (.O (d[30]), .CI (nx62012z1), .LI (nx62012z2)) ;
    XORCY xorcy_31 (.O (d[31]), .CI (nx18600z1), .LI (a[31])) ;
    MUXCY muxcy_0 (.O (nx8474z1), .CI (nx8473z1), .DI (nx8473z2), .S (nx8473z3)
          ) ;
    MUXCY muxcy_1 (.O (nx8475z1), .CI (nx8474z1), .DI (nx8473z2), .S (nx8474z2)
          ) ;
    MUXCY muxcy_2 (.O (nx8476z1), .CI (nx8475z1), .DI (nx8473z2), .S (nx8475z2)
          ) ;
    MUXCY muxcy_3 (.O (nx8477z1), .CI (nx8476z1), .DI (nx8473z2), .S (nx8476z2)
          ) ;
    MUXCY muxcy_4 (.O (nx8478z1), .CI (nx8477z1), .DI (nx8473z2), .S (nx8477z2)
          ) ;
    MUXCY muxcy_5 (.O (nx8479z1), .CI (nx8478z1), .DI (nx8473z2), .S (nx8478z2)
          ) ;
    MUXCY muxcy_6 (.O (nx8480z1), .CI (nx8479z1), .DI (nx8473z2), .S (nx8479z2)
          ) ;
    MUXCY muxcy_7 (.O (nx8481z1), .CI (nx8480z1), .DI (nx8473z2), .S (nx8480z2)
          ) ;
    MUXCY muxcy_8 (.O (nx8482z1), .CI (nx8481z1), .DI (nx8473z2), .S (nx8481z2)
          ) ;
    MUXCY muxcy_9 (.O (nx60018z1), .CI (nx8482z1), .DI (nx8473z2), .S (nx8482z2)
          ) ;
    MUXCY muxcy_10 (.O (nx60019z1), .CI (nx60018z1), .DI (nx8473z2), .S (
          nx60018z2)) ;
    MUXCY muxcy_11 (.O (nx60020z1), .CI (nx60019z1), .DI (nx8473z2), .S (
          nx60019z2)) ;
    MUXCY muxcy_12 (.O (nx60021z1), .CI (nx60020z1), .DI (nx8473z2), .S (
          nx60020z2)) ;
    MUXCY muxcy_13 (.O (nx60022z1), .CI (nx60021z1), .DI (nx8473z2), .S (
          nx60021z2)) ;
    MUXCY muxcy_14 (.O (nx60023z1), .CI (nx60022z1), .DI (nx8473z2), .S (
          nx60022z2)) ;
    MUXCY muxcy_15 (.O (nx60024z1), .CI (nx60023z1), .DI (nx8473z2), .S (
          nx60023z2)) ;
    MUXCY muxcy_16 (.O (nx60025z1), .CI (nx60024z1), .DI (nx8473z2), .S (
          nx60024z2)) ;
    MUXCY muxcy_17 (.O (nx60026z1), .CI (nx60025z1), .DI (nx8473z2), .S (
          nx60025z2)) ;
    MUXCY muxcy_18 (.O (nx60027z1), .CI (nx60026z1), .DI (nx8473z2), .S (
          nx60026z2)) ;
    MUXCY muxcy_19 (.O (nx61015z1), .CI (nx60027z1), .DI (nx8473z2), .S (
          nx60027z2)) ;
    MUXCY muxcy_20 (.O (nx61016z1), .CI (nx61015z1), .DI (nx8473z2), .S (
          nx61015z2)) ;
    MUXCY muxcy_21 (.O (nx61017z1), .CI (nx61016z1), .DI (nx8473z2), .S (
          nx61016z2)) ;
    MUXCY muxcy_22 (.O (nx61018z1), .CI (nx61017z1), .DI (nx8473z2), .S (
          nx61017z2)) ;
    MUXCY muxcy_23 (.O (nx61019z1), .CI (nx61018z1), .DI (nx8473z2), .S (
          nx61018z2)) ;
    MUXCY muxcy_24 (.O (nx61020z1), .CI (nx61019z1), .DI (nx8473z2), .S (
          nx61019z2)) ;
    MUXCY muxcy_25 (.O (nx61021z1), .CI (nx61020z1), .DI (nx8473z2), .S (
          nx61020z2)) ;
    MUXCY muxcy_26 (.O (nx61022z1), .CI (nx61021z1), .DI (nx8473z2), .S (
          nx61021z2)) ;
    MUXCY muxcy_27 (.O (nx61023z1), .CI (nx61022z1), .DI (nx8473z2), .S (
          nx61022z2)) ;
    MUXCY muxcy_28 (.O (nx61024z1), .CI (nx61023z1), .DI (nx8473z2), .S (
          nx61023z2)) ;
    MUXCY muxcy_29 (.O (nx62012z1), .CI (nx61024z1), .DI (nx8473z2), .S (
          nx61024z2)) ;
    MUXCY muxcy_30 (.O (nx18600z1), .CI (nx62012z1), .DI (nx8473z2), .S (
          nx62012z2)) ;
    LUT3 ix62012z1498 (.O (nx62012z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(21)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(30)  )) ;
         defparam ix62012z1498.INIT = 8'hB8;
    LUT3 ix61024z1498 (.O (nx61024z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(20)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(29)  )) ;
         defparam ix61024z1498.INIT = 8'hB8;
    LUT3 ix61023z1498 (.O (nx61023z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(19)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(28)  )) ;
         defparam ix61023z1498.INIT = 8'hB8;
    LUT3 ix61022z1498 (.O (nx61022z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(18)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(27)  )) ;
         defparam ix61022z1498.INIT = 8'hB8;
    LUT3 ix61021z1498 (.O (nx61021z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(17)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(26)  )) ;
         defparam ix61021z1498.INIT = 8'hB8;
    LUT3 ix61020z1498 (.O (nx61020z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(16)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(25)  )) ;
         defparam ix61020z1498.INIT = 8'hB8;
    LUT3 ix61019z1498 (.O (nx61019z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(15)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(24)  )) ;
         defparam ix61019z1498.INIT = 8'hB8;
    LUT3 ix61018z1498 (.O (nx61018z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(14)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(23)  )) ;
         defparam ix61018z1498.INIT = 8'hB8;
    LUT3 ix61017z1498 (.O (nx61017z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(13)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(22)  )) ;
         defparam ix61017z1498.INIT = 8'hB8;
    LUT3 ix61016z1498 (.O (nx61016z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(12)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(21)  )) ;
         defparam ix61016z1498.INIT = 8'hB8;
    LUT3 ix61015z1498 (.O (nx61015z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(11)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(20)  )) ;
         defparam ix61015z1498.INIT = 8'hB8;
    LUT3 ix60027z1498 (.O (nx60027z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(10)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(19)  )) ;
         defparam ix60027z1498.INIT = 8'hB8;
    LUT3 ix60026z1498 (.O (nx60026z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(9)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(18)  )) ;
         defparam ix60026z1498.INIT = 8'hB8;
    LUT3 ix60025z1498 (.O (nx60025z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(8)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(17)  )) ;
         defparam ix60025z1498.INIT = 8'hB8;
    LUT3 ix60024z1498 (.O (nx60024z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(7)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(16)  )) ;
         defparam ix60024z1498.INIT = 8'hB8;
    LUT3 ix60023z1498 (.O (nx60023z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(6)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(15)  )) ;
         defparam ix60023z1498.INIT = 8'hB8;
    LUT3 ix60022z1498 (.O (nx60022z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(5)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(14)  )) ;
         defparam ix60022z1498.INIT = 8'hB8;
    LUT3 ix60021z1498 (.O (nx60021z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(4)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(13)  )) ;
         defparam ix60021z1498.INIT = 8'hB8;
    LUT3 ix60020z1498 (.O (nx60020z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(3)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(12)  )) ;
         defparam ix60020z1498.INIT = 8'hB8;
    LUT3 ix60019z1498 (.O (nx60019z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(2)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(11)  )) ;
         defparam ix60019z1498.INIT = 8'hB8;
    LUT3 ix60018z1498 (.O (nx60018z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(1)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(10)  )) ;
         defparam ix60018z1498.INIT = 8'hB8;
    LUT3 ix8482z1498 (.O (nx8482z2), .I0 (
         \p_reconstruction_error_for_for_c_sva_31_9_2(0)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (
         \p_reconstruction_error_for_l_sva_3(9)  )) ;
         defparam ix8482z1498.INIT = 8'hB8;
    LUT3 ix8481z1540 (.O (nx8481z2), .I0 (
         \p_reconstruction_error_for_l_sva_3(8)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2488)) ;
         defparam ix8481z1540.INIT = 8'hE2;
    LUT3 ix8480z1540 (.O (nx8480z2), .I0 (
         \p_reconstruction_error_for_l_sva_3(7)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2489)) ;
         defparam ix8480z1540.INIT = 8'hE2;
    LUT3 ix8479z1540 (.O (nx8479z2), .I0 (
         \p_reconstruction_error_for_l_sva_3(6)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2490)) ;
         defparam ix8479z1540.INIT = 8'hE2;
    LUT3 ix8478z1540 (.O (nx8478z2), .I0 (
         \p_reconstruction_error_for_l_sva_3(5)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2491)) ;
         defparam ix8478z1540.INIT = 8'hE2;
    LUT3 ix8477z1540 (.O (nx8477z2), .I0 (
         \p_reconstruction_error_for_l_sva_3(4)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2492)) ;
         defparam ix8477z1540.INIT = 8'hE2;
    LUT3 ix8476z1540 (.O (nx8476z2), .I0 (
         \p_reconstruction_error_for_l_sva_3(3)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2493)) ;
         defparam ix8476z1540.INIT = 8'hE2;
    LUT3 ix8475z1540 (.O (nx8475z2), .I0 (
         \p_reconstruction_error_for_l_sva_3(2)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2494)) ;
         defparam ix8475z1540.INIT = 8'hE2;
    LUT3 ix8474z1540 (.O (nx8474z2), .I0 (
         \p_reconstruction_error_for_l_sva_3(1)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2495)) ;
         defparam ix8474z1540.INIT = 8'hE2;
    LUT3 ix8473z1542 (.O (nx8473z3), .I0 (
         \p_reconstruction_error_for_l_sva_3(0)  ), .I1 (
         \p_for_for_mux1h_2_nl(1)  ), .I2 (px2496)) ;
         defparam ix8473z1542.INIT = 8'hE2;
endmodule

